`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W3GQ2cphRiNtOf4YSkhfjXNAbfB9igv+tZQdLj7Ui09OGMPat8fP3KASw2maWD29ouVKkKLvG6Vr
91PR0qdglw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gZ9c7DiEYAEVqYa/yMMLOD0vExaRRYpjctkFZRuVbqn0sVY9GTNCExEYOaa4seaaj8EXXpIb2S/0
YqQqAHPjiPoIBLmcVGY8d+fbMl4LsUaWFwbNMjyrZTI8TA4g27x5ofBuNx601IcCfx/3yqJvm8wL
AJLbyzpD3cQVSryQXEU=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nbujIDXvFS5VIX6eTJ4NmsFeZbfoQqCXaDKqXGs38PRuDJs0mDuQN5HYpGeqQSnsxcv4AGRP7CKl
8aB3r4JmPRzogWegHwLChYILL9J6B2GQflyW3s9Bq3R+YRWmtoT/cJj6X7L452A+zzBVFpmACzU9
aRGmz+VCq3th2ki7pRQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BYIxzELlFwptNNYbqLbUIG0VOw572GbHRl+zq1MRbtEO6coJqDuh58U8ZH5o+Oh3B2lZo3kPlcyj
9QqGtpoVFLBWAIWxkuLZTbejClImJx0NpZOsWWYqcnNEnD7vz1srqKcNeRd3jKI8MnBUgKk3jrLo
HQdiDyaKdXQ7lB9TcpUiWXER6urMzKPvkj35NcqJOfcf2NgQuPnC1lVABj/rvrCXlNhZ5isjSwSA
Jts40np3vuLLp5Rp17ZZpGAPDy83AZcF93Yu013ZjgKYVG8uVyYoNTvR7h85Vp7oTslRZ3oj4OOf
/eUz3V/KjQ8FdgHzS9damMZrvYTKaNpRNr+X6w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FRRAnnwjSzbsDwJz9n1ruM4+OWqYgO2yiSUwMwj6JVaMDzoWgBNMXP+5hci9QJdJplEEhDS+KHhF
Kq8X8cm+aIE7/ibWb9CDHwXprT7tYnp+6A8dBMNk/W5Spp4+sk3rlPirboBaJB41KYyubDCxrgXf
3DyusmRICyAq60hF7IOHjGOoqO7oGOMzgt6XYLa53nYIXJdQQRvbetQt0watabv/dNht8FQtXj8v
O1laGsl1kMeGcvRt8tKIpbQMnq8hubZJE5g62Ou3E6EJMrEHMW8Nm5luPQmo/b4i87Xh6zJyzcbj
W2jHb2quXeYh8qhu6qc07re7wuVY9X0SKtMPhA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GeJIhuD4RCTO/yzX26HYXpttHs/SUokwH91LoXenqWkWNG1+n61IO+vs+kb8GX2HjPVOVwg1ulFj
IxdoBLOgijmatLNlrp/sSuWzjRZNKD1lTdzd/6/8f1OzKFfaJ6dFWC653yEWEzUTPIYX36fqTxdw
t/whcIUWfGut/EzGau5GyITBD952jdSgI/aPpY9q+sKb/j9qD0xMxwxP30QXJiS1Q1R5j6rYat+K
dXByw8Bofn8M5/RF2kduY4YZNwawvjguR/1gvymUjEmG2u6RWt/OkMSB+2almzIet+tKuoxo4VH1
VjBpWVmnJ3So4e+Y6OVeZEC+DeRyQQGZYKqvTA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 648640)
`protect data_block
1ZgoZ8xrYuPlq4syMA9wBNUTkYxx69qNOPy/nj3HiSGkaCgd16Po5HrIH3V8LyJKEY+ydAUqKzkE
BX8ip7MEPjkS2h6KkNzoiRvNjcW0Okj4eqtFVcZo3QabNzFc4yaEoWrIlf3eqSD9t/sUqzhBnvm9
qvoF8cGtn4IRYTPYQnFBuU3/qptxmB96V+pkzqevTK+SFgkjG1FqqiCd/Dx/loAaHcEQazRTS9xf
n1HNmOSdUoo9X7Y+H3ZT2i/dn+N6vswV5lLTklDtKyQ98MRjeKTa5yxBdufMuWnDOcmmcA1Cdq/M
nMOEUYPb/Ab+eFr/T3uQIVWFUQEOf4NoiXTlPerpO07kLM2EIoNj+rc/HNS7xBNEatImSmdTzazg
pYyqg5nnMB8zVx0PTVlId9b+M76stR7fnU/iAEscccMtKzADvi1THi0kQZEAJeqyO1f2mehW4W2r
LBZfSt0Z3xSGY0yFKpwfZgr5fK5RO3PBAruRHfDKlYwfhwGSFG+hvOOfC7aXF1Cxu2dPC2zb0P0u
NRlQR/eJZYGgJcBHHKORIYhh/jIQPb30nbFK6/g5g94jFJDOUJtfN6o6ymf74Sout2jP1gV6TU+X
ZwtixjwjdCR41doJqwXLyCc++FqezYaBhY4wEykTZvdUexF1k7tjfTQystc9iNYHHT7nrt3aC5JN
vADau3xzVDSE0HoCZrv3fIlngnwxjOPjod8PE/5MRmL6WguRCgEHDKzYZwO7k9owcSX0D6XRMPDZ
F3PMO+CSRTyy4HsSyqCdCxYEk/D++XEzPswUiQWAZk7YoTas14U58NmVjAm0uXuM2ilZ+SuCB7DW
z6BOxExGD+Bbtt8K0S5rppoGO0JFvMZAUd1pkXV7niYHiZRMPGcXBsC8eqi4fysBzi16MuNwUaGD
BI0jurRCrFU1VTQbq9bjkytbEuSShTq59iYvyqrf67TZGkwtQ+aO1QBSDuZzkZbflGuPe8RDU67g
4G1lA3iSRIhRSTJHyTvl8sMk0iB+/buJ7BXttIeloMtNPGE2+jo/xwQh2oRLdM885pmI7X0r/EjE
vaABDTt1Ih+u9aCPB5kBarNZoLRp1A22fJDY8gNW4LsaNIWwcjV2h36JzwiN4dvFoSY+8BugPqFo
lX718giB6uK5p7vMoBpd34UYvrgxU13QC0DiS5LVZCEj0I4qTXJxI73FdfCJdvKPCInhUGOTxpmH
Pvi2QHaIJBUqu+snP4mI4YVIcvt5DoWrevM9Qzqz+ej3D851GwjZHdhfLAH7V14QQHFa/l5o/RK+
nhe4+Wbb8s/SHt/H35wzHl/3l2vwjgQGi8e139/lJR7r1laWWlciVV4EUzaUXSjmOk08aTVt+I8+
T5mTKlB0s4KdyVrinKjTc0RMkfMkqARmlpkwbph86Uyjg+moERUclTz4H8nxGiMiqZsunE9I2D//
MvhyaZSZGTRfQkqnsBslKoMRxTdRQAZKT9hDVdu9lDH90U0R4IOGOHRBGfeMFTQZHEB3OM1Bwdaa
E9tQ7ewuH8IYW0tpG8HBrq9ultlyfrnmTQdb8wcvo65HeoC90VfgFXtLGe3qs7bRUJ+VKBU2y5fK
TWcu3ew3SIyG61mSKOooYH8LBL2J43xjeNHP3mr+elcbizVmN6MqUD/KJ/ec3o4g8g2XI2rzZ4EK
6pJ6s3ROTJ7hfu3TcleeRvSYnUPVHOXbppCQrUbaSbdm/5XXEdbqvBKZ3VbVU0W+vbboj8zJ4cwD
r98t3wBo2g+Vur+xEZJhgKbllPdxI5UfVxHH+PM9LT4Hy6ibUHdU8c3oA7H57FC+bT2C8gYO+9Ps
VIjFzdx1OBG/zz2CNf+DZsHBWKLPZORqbuc1Lw0qUKDoBjX+AaMMgC3bFAPj6rb0bYt+uVmx8jyh
+aBUEXg0QctPdJfH5umTHT6+FyOc3+kL2X/JoB2o3q+ZIC67Q1L1wRahH+MkLFUVY9z5SFU2iLFY
gG0qSLSLoq11DslbFcqufImnIYj9kR6BzrDP2vxcrDC2eCx5yPi2H4oVpnDAwNPzUMLTZD6lgrwi
oz5wc3PlmORh/eiZJGuwovktWNnyO+rAsLNbcyP9LOs6Lbikfo9jC32bJ/XtrS6lpKKGjv1QVPkS
10gzYJh+wLYiW1OrA/TpQcGGUK0VqT1o/R03Btea25USFCI33eee1XJmNjXHtQqIi2oB4eKbgdJZ
5qxveZwRU+hgOOdaJXZf4W+j2MXoRTZoCOvwSDRdUGC4Zw2RThi+Y4S/5tGVwQapaw0xi02/QPgA
NNyNGex0dFWprakgRytGe9vTn0XWmjclaF+WnuLlOYE7DoSc7A0W2HVkFgAgT/CGxaQqchkIIl38
mkR8RDZwv5ZX30XZAJ3LjuYD92tR1quWR+YzAfbN5UQtkH8QINCAIjqREx/MiB9bKwgyK4VMS44s
NgCmT7AI9FBtx9YbY2Nggi8aNk/gYzfln7t08DjYH7ru0GtWdELIiDSbYcNxBxKYFZ/JlqlSF96M
yAYh8KkQmdBrDJEUYu/lx855RdDQ3VbjBOf93sP1VXO+p5f1oYtLzgxu8eSLZublgjzsTfXzZdaa
2xCYArrkL/GQT1ED+JivfBBVppWnzy3yFN50VfmTX4PjWWyPQr8PcNSJSVXkRVbAqdLmNV6a4Nke
Ulme1tOg5o/fFvf6QEx/tztvwPDUxyHvtZza73M1HuJl+Tgy9c64TNZBxPnOM5LXocYhD5V48H3M
iFFtSwIDQSj4ARh0z77xLNKEBibu9152xcZs397aPnv6yU01lDCDAyTX+oPvX/qJAseKBnSSCFSV
LVbhTbVsLmXlsS8A5CZqa+0vFiLZk58nlhqPDW/+0UCszcxoR6Coqz7kLCitVTHzMX38Tiv7jhVw
Z+oAAz6ofKrYNiwOS2feoHfOxl92ZYTBy8r8gpXTRy0SXIHtjXpeyn7r1Zl4UZwIE5tCeTlVXoPr
SBtFFuWWjvegDF6k8ny8I6iX5jdltz7COk50ZyJiMKVQzXoqaw8Y1KiZIE2OgOc8WDLs0rqe3AEO
usVIRwUwPLXMtMRnPWzDmW//ZcMcZb7KmBFT+vc2GfIB0EaIskQhhQbINfBOfYGLRo6M3mZSJ7Q6
aBFJSwvEGfLUREBHND6BqqZqGhIZM6Fwn94lF9EMPCbQ/3kce6ozKYTxvSVey38DlAbUJp2UGtlu
axBdYEP/ve/CCqfygrBz919IMMnI9IZFr26j0btRfQScBvXhn7iumBZPHNPIZHZ3y5UO3Ou3hiN7
mguWQLrtGpyOD7163M7wfp5qeCiZVyxfb3gLWWi46h9Ow4DmMUkFdzBxXRajF/y4yPxHjLxVsyNf
LjZCJCeA2pBSdAEiA8w6oS3i0poac+0SkuwdNBy3uZH5q/8DJiPL8/9Wz3pgsWGiU3Ci1Wk15y0t
qExWCdRQZtBSde5tjHaF1ZjhzpRDxgSPUlwYuHybioUhuAnAPWuIMphsDtn2u9wKYmIz9g2LKQI8
l0zJvc2k9GljjMfrNaYbuKpeVwROtpIEKp8tSTgl2Y+mD6ZRRqwiTK1EQitQq++QBcpkEHe8Ucs0
8FAYVTh8l7LieUQzs7S7yI4noY7jdH/5yI6E1MzLooN06RBB6TIM8imwvdIYzFUiOz9LDHSQ1ffW
VV6Wx00634TV6pPihsB662U6d9Y5WSSc413VuiFq0vrY7DsYDa0JBKkvDOTVtcKHOEl8Rxv+Th21
PNlJE6lPDyMZNBHmj1+YFYzhqnW+BD3YTKbjsjEWeItQqJcOe6qVgOhR0W/xwh85s0N6n8nLOEYT
pbYuLNymABPUMw83HOtKigiM+QdmUMPyIdj1yzk3kz2EOMEAW2kHaU/cyrE8m2pPuME2qt0DpJCX
zKHXeq7p6zcmDcJ+MlED5MTtMnCvLN1ISIQRk5TGMtmvMNUAIKZQrhrBMl6tGZsYNH/dq2C2k2lC
6iPuw021mnRB3dBhKk4DKd+v+AKfs1V4GlB75NwdynuyjhnbxEtCV2YHuZoaCaIDMCbk6GjUKmsF
IolBanw7Nm4B8g1SZWajsIxHSRG8LqCQt2qcYzGYc3YSstIrI0sfOLj5TUv86ZYdWYEvttkrYndu
/nFh7pftI5KT6sH0iaCcwq08OG7G+RhlHS0VXr4cqzPyxe1gnUghINwgQHNbJ3Rz4GXQUNhkdRIG
7ElTLuFCAkD4M0Sk8k+jGvU+4cUV0wadMPncBfYGoK4Lbq5UBKTnXcgpyNckIgbYm0/8QaxAI5V4
reOpFpU71hDZZGiFspVQFt9/kZEi1UUftfM450HUZQjMo90eLDDP0CVM5z8a6unRrzrGVBciASy0
2yhlo4z8Wz/YTbJ43or1vDzW2qbWJxqY4jg+ZqYxEPrBiYpCxS5kCgholMhQe/w/X+jcu//+h99Q
iNEO295L9B3WOWg7Bs/WeyLxj7t6l1YoUx/0QifPJTgVLpept7zsMJkbtn5AL41Q+N1k4xRvWsRe
O4p1GCPwAYG2tXXkWWMMYq3NrvaZ/IOClvBqiXcSJpHx/GEqnkGS6/bB5hKJRu1yMrAxZT2fXDgK
omzSefkDYBw09bsSmRJOgm0JVzbO4RqUwXFVkbR5NY1862Th0GF+7RODkK/jfJo99lJMj/TdBna/
E+dHKgo88MDe9kqI5ESTdaqm7NSiWqZ7HOrEKYRSllf2dFoFkwl4VzpEgSBTOYZvndwWX1G+DTmU
h2nP5VfPU9WKmnHpV7ZEg7JT1wdK8ZbAIl8m5MxlhMjW905+wy/QbeIgnuCNQB7Mke50E3w2rTkd
lfU7+dQgt6gmO80N0WHeLWPsa/eoJeBp9FxzhBKPzSnPBc0vboDvN4w9ifx2xJNqzN266cSiK/ol
5pRQ+UEmK7raMF+exLMZlQn0tKkQwRxSaeJNWDle5vu1t2nGAeX2apxtoo5ayVJMjWJ0QucFEG0B
7wXl4MXReqpWZpvK43YcMW48n0K4yDYWm+x1QUtmp1ibM2t8wXpcVSuuvP3gFsUMetdufHcLotwW
srRALbXDTFaHGQ4o65ZfKNU8h4PRSQeR+p9wRVNFQy96j3WsLMP0AcmSYbgHb7P79gfFbLs+EVbG
DLIKh9vS0ADh1kIKwdNh/9hW/P+zJ9/1fwaklV/7zdKCk97Bce6rYWek+coacC8Z0cc6uRMWt4JQ
PTTTqVdtH3efq2k45YwXC7mqTdJSax9i64vYyuOrREp8H2TlbitDT207vhw24nCZa4KAowIykRkK
rLyn1fQvE9gmIvTjIeZ0j+fAurdpCWnpeXZ29/61Kymxo36S2yAY1JY4CIATbf/KQVLyUO9K/faH
IZb0zDdlMiN6QJ5jzN4vuRkZjWopsoxRO5GUzZK1z0d7qoWM9VIwzArGeAX2x7MSQGnCgRX5VBGr
8fMxL4L0dzvfKZJ2n+nE3fe9UjvwXhLKItsyCbjMZTL6lb9cQB5hUqggvXQVKuk9ySv2JB8tUDRr
R7F4MxxmIGM+wCs25bereXwucV3aAmAWas52REFtEERvdwlzCpdQrMctyGi1jj7V/MbWMCOQoRJf
BtOyFGcSEvsHWyrNt0u34pge2iPe5MxJtI86SsCPNhPf51El2Htf7J4myMwKad77hrlwEk+XL7K/
rvNiIBSSJX/rTPyLP/626Po7cQbH7dRPCs1/LSOaNnaEM87LiXXwLy5tuVeECWltrsKrAXoGkO6s
gcvPRHG776I+rF1ou8fetL0mNtaaLd5SwHAOVKFaNmRVJS8bozV8w8NBh407ZaXVwKYfRiKsfSsa
esYwbSoQApI0BgaINKOhvOlbuF9wkzJF0RRRc5fETvfbQd++zkliR+pEoUG5LffgPzsC8+u76Ra4
02haZIae9/8iv6agIfRPB276kHwP1j4bWMqjRgpYgCb+QonqOYfX79UOPWgzrZzaHI6H2SwCCwG6
CNhQIvMpRTacq5HnVvuZTkbO+CtDtQQv0Z11GNa+VDc/J4HYqERk/9nx1nbDVYtO5tvCz4Y0gnn0
/5ilJ3e+pubYVIaLKoVlCD8JR0y/SUwxHEyrkcEfWUBvC7Sv4SMGh8RroFNrRIcAkbudjZHXA0mK
U6xqFZzHbMZig6uf36gTZ25x6mCxo811WRa3Lsu6CkX6/C6dRcGFnEz6kIBCNFgu/DOisiHzzho/
umIw+L9JhMJaNqiR+bVR70KGKIZcuTPjRMHSvy42ipjxHNTpIke7IfWm1Y18XQ/LBDnE5J1S3V+9
0pAUFhXnzboXSJOXXOBGeEe4oJa21yaraGvG/pd/C/ggwSGSFUd0g4J1Xdm/TRWGV6eYK9jztQnE
nSevijUbGMvNRMvIXmlAnzaQgH0bsXLfYc7pt8mMNWtpOL3QTBpKmv7rHmV65EbHXa6IrXAxydFO
tYCxlpMR0ncwJ5TP3qSWZ3NT+a1ZpDDNzLkGLl+SKXsJBVrL6zAqStPtsqJw2vuMFrSU/+0PUpLL
4PcA7fqO0WkLSp8FZQa3IGFcAQ1UavRCfT/mdwgKrpC1mVe92aUv5bccIcvtU342f6gNamOYzHKd
rxvx/acX548Sho1Y5R7bjxQn6gyidHXUNo2KhV7yDONO3rHXH4j1CJV9gNU3vXa1Ad4yWFCQRmRG
9TuOJAQPqRRbEKNadLcu+Z1JWxLqYsQ/Epnj2X8e5qtK/U2LJ8uRVC4UTjdamj4siXpjSK4gaDAs
Q25XgETajNR/WjW9s8NqERrCDUUKvairACyx1FCBLxzBJFa8bOMPjkp8HsOfDgr24M94RzrIfHLC
Ov1cIe12FNap3/AzXEzqjqFsK6ck25FhAYXokVzH8tufVx3Q4etukbgyZIm7XPAuHF0IObbuxXgh
l1NdO32cr63aOxknDjUml8aDpM8x6v+w8oFh0dM0LGWh1M5fFc672r1jYrJt5HUoqZvNoED+9URV
lDVJCk5mpd0TpMWogDtR8NNbr2yiSKHiia3mswZ4zVuyiyfDWOHzFaOxk26Ud5Hd2hvvZ6z7752i
8cdVaYtkykFNCh2xNTnr2vNyuVcnr/mRaSFnOeg6qsDnig4rOYJBsXBRfcBG+2L+0Wf6dS1TJfXA
a7fDqBd/u1cYpGrvkwQ/25+sNoQ8mFBQ2cowVb11xf4ZrkhtPHGeNmvoAh/1rT9ThukMe9xOFd3v
AxT80AQNYvSMcRGdtjd5p/in2IjBYN0tgqPBwYi+VONdX+QpSF0qUHKpCOTwrPJDmUNztBxiz7pQ
zCrcLEMnYsEE8QK72KM7YdODKGZtKrZ/wOJ5GTzKjEVjBpkbi5BLI0d3QKnV0vk88gPFbiEsNVRf
2Tk3UGaeXefATJn8sShW40Rs969X6J3yNEJLdWMbe0WcOUymG6pTCxNXv1JanX8eIYLjRE1xwcqP
W+GX6Jizf7zScwkKraWv62Upqt366P7eUuGLBTvFKrAffdarjrCBTEQQ6OpXEXI4EvWz9H8CmDDZ
1hs0ud8mGdBIL+J6dYQQhZqVzmb3MrAMKt1l/gnDAqgVd8zpqF7k49r+GN2nBOCfHPKCUXsIvPIU
hRom5uCkq0imCnnMEYQ7iYnsOud5m/qag3eDiN/jiBsdg89FZ1DNdsgXDWGunPU+67hFD00XRiWv
ZRDqjwkjwMS3PfeDjP57Hz5mwMbmtbcis3OTEN3R/BFsS/aJB73haC/x2leI9GIVf4qvodacN+3w
Qide01O2F/IxuMrX22nbNaXJIqiaV0SZwOGg3WYZrnXDlMMEgxDK3SOvWpz1PObc5iQ4bN5xhxxw
D3I+z2knyG1AbNGlad7wsyDQwemol2wt3MeE5lnHSJjcJr567mvP0hGiT31oeF7ECKW/+FiJACmc
bl8nCnUbq6cza6DVXD+PLORqw9OqCr86NUeJzRpBxYM9jA9K9VUP/wQwypirfnYYBgH/ZkrN4kM/
3Tcp9GAtJRHUD8ZKkO4AL3iFtC5Nr+YzWaxyWMYC7JbTV3q+1vbIuBmBemurfGqeVfjm6LTz1MNG
wLZTqVN2ORp+gg+c3yiHG0VC0VRczA8aLK5O8vKp4FBdyQy7QGJjyFn7h2gcjVlNXUkQzaK4WiyF
AeD7xuPmyWtmURiFFOV2XsyrabOuB3uPEmjFYHAWPv7KLYF1d7SS44iJXdie7CEa18wDewsqoWvC
xG2cCrA37tCcepL9BO6aIrvTGmbCQsFZWy/GSd2q690iDOYfWbme8fmmSSFoYYO+rRo7DZHCK3xy
mTuuKMJaUQSVpHsMNmiVMns4bowB0ICQ6qydnxfY4IF2Ya0KCAHNlI2KruJzt7kFK05MXgdI0UqT
AMVsNw+tkm+M+ifkb8Yr9zpmrLfO3KvB4fiXa+q138h2Fj0fnmEdgBMnOBDFcXsuomKSYoVS6vMV
RK1koVWozglfF51y/yW4Wg1GyAMrov8SeYHRFcgO01kWfojG5IL85eyODf493JDsDwB3vzakzCoh
dENGwoiY/z5S9vsUfuY4Cj4L7ikxuR0mvCTBv+Ha4mz0jGmIXsPx4BHGq14zLJ+1KY6WU4bT4g1g
YvwE+jOCn3RaqaKB39zwohPnd6iqQAeH3t7OOHr3w7TiGey1Bma944e+bzJkWoSsA/W6Ma72/wFu
otUDNiSz/Qt+PV3XRgrzBMfGwMyIR4W2ycp+LSZLgi/jFTHqcTOF6HoAlgWCS0q7Zj2SDIG3CHKk
RORI2y/cibYynV2WmtSrhYj2wSH8j4ZH867cFQ0fTfNI/hP53bACIiBjxzab8T5l9raDcWFXUck2
9Sj/pRaY6GvR0P5yHlu5LlpizfZXlF9hv/B7pwTNeEx1fZO1MUOTmztNbUOZR0YQbysLAvtHo8DC
qWGBO/n5ML+J/PBcLtKw08s0ByXFuudqIVeX4ERBs5q2R+vPvGq1D7vZoHeh3X17Z55m0Wx/eIB8
JwZUToKv/DthVodMk/+8ZofHXyXt7JV/mL01P3S0K5bBTxWC4xOVQci+dKDT3yeG6Gn2EFr7tvd8
gltO+ILrnxBNngZOqpg9VqghYWb/oQ5jg2Zwsyhsg6ooheR+UzycYUQOmGVdykGjBvyVsdWR1YIU
6kJKxqxcb+wO0fk3zTeLbNesiHcqeL48DmORG2YM5pGeWTxJjQikwedzmWyU0QgL6eabHpS8xJfX
G5czo3SzNDaIG5HMoqPzI3yHz/56nPZJMr4L44h0lVSh1lSJgSTcZ/38yDU22fRp2fmMxF0tJs4O
8+qqNwxSC2TcyS6FUSa8ASVHUe2V6mEyCOhEwM+NvhbrKhPD4eji74FQ15X7yBYbzGx6YXd1jnri
TBKwpw/YoIPScpNG2u3siXrkCktW5Pbs5fRCQs7JJQJB/Hr5s8gMfeE29fJMHVL0fnlonLlIgV1+
pz0QaE5y4leWNNpE0LFQlrI4xYdvkzJElhv1kuTXq9rNaBUW90Z5h5vdmIQDh9qkK20N5wTkgH8P
7UOiofUNyH/kjrnQ5rxtHAMyack9jeJvOzv/KF0jPtBeRqRph+N7hkHRhRPUerdzG9C5rZwea/cS
EPC1drWsh73fMkvevwC9ilil0HSfLGav1f0BR41ASMsB/iQDEJY3Kk2gtcuu/FkMtidwYJRaYncf
mG1zoAThwes2lGlQDKI5ah8+CB8zCIjnSZAkc06NDBFWHi8WD8wdgh3BJE1uUBFmxWZRSIWLI+XC
ioyPCDfnBIvfEqlOVN5W7BaCUY5mEU8n/bZg/29FwXhx1aP9Z4ovbT2uZmEJZZTyAUT68hss1IWz
X6eAbo34+W0ba1L1qktqc+3MaILt3faAiRFWHDdXnSp4OR+WagSC6/FNRgItWA+xPzE+ASbX4JLe
+ppX7R5PFEJYi+8+T6C8dHsGxoryqQER2MIhXAiCCWnRwgO/iOFoqM6H8T5YWIkc6XqWbj1N1bLw
EuYF8FX+EsulZrwXH2H3uk6RTUVhGVAUsVMkOE7E5suzvZVnBo8Ta+TD0a92G69j+6Q0XHcq09Ou
+sj/z8nn4zbrU8ZiSoHubAr3HNXGt4AWpp5kNgWMrAJKEYNGdSoZME8NxlzpBQ3JcWbqDeGkNYgw
d2tZAx+siP7fUAYAJksSvl0LuemyzZ1wVvSAhkHyfgMyomGoq+PVkueT0gH7W0a07d5+lpUDOe2J
BfB+Z8xPumQZMXtFty7s8YuelTFoQMAs34HDokacovFjDq12mm9w27quIK7aJx3kMHyNqzLOEWtp
9qwsbfbd0fKWNdrFwCdPxumsU+k4bKCTFopwMqq0yEVzYDt+RwEgVLFSw5n6AVbIGUj6AqkhipAZ
ZhviSQkkdGjkheBlyHLqfKs22JFfllqzRiEbkswb5TA1HGuPFVxQXmTiv77f9tkzvLtX/K6TopWT
w3gjaibIpuFgoTtxMTYGRCgOe9RxWxWSgB4H2HzVBNxLMojdvANS1xND2BKogxMh8tbyDopIyuyB
mCmPanQ//g4FPJDPXbz8SKMZABI/vhaj/mR21mQijUmQ+1nhFUy81OqSR/Xv6WkYCA6NBwbwQBXu
/PEMCYBrOzauQ+xGzu/8aVrmgypsPtXUhAxWSCm2i8MtSDcGZ8l8lNIsbhG/51fzjoNzIXmMs2JP
cYM76seUqBUvaqTNauFd5jbO9OoSMSizRWs5n/As38JMxEG4EOWE9NikKpfZhAApfn6OQVP4J1pV
tyf9BFIqyXK8EHFuB/yt/IgRnA53tFakmlA4O0CYxQsbzKAyZ77/LRh5yHra4nyZ12l0oprFxInG
Nc0Sg+x28OY+BHQltUaL3sQq1PTp3YTmnVu+ofxM2l/fMUR48BTXm3FPPqZh6EI4nDcExEyKj1O1
B0v0/chiqGUCXzLGFz6l9nwmPxryIOGAI4JtWZ2HnTyqZUe7B7OQ59Pm6oTMha7FshA62nrVlyuP
asFNkqcSQZTrS7i+JUeuQI5rIJ12AqdqwJU6tEiOcKuYk6KFI1xnvPRMWLuYTGCB6ElLyp7Ns4Pk
KtW91bQQ41fcOCXM6wJJCPjB4zgbdg3S2IoD7KoJJyry5b/ha49PE5Ju/Ckh7Wo9vc+t/EwbWfoT
IQ9g5WWWCMkEjcdoao5bY3/HDukQlJSrJ+wykVC+BBsGnXU+28GYOepX5x6xBl+sc2HPz9KgxDJ8
zWesjkWrjWVcLTOQIty7D0P1l5BICDowCUhvLahOl4IUTY2uhy4NLQLzfYiQc7WYLJhvOfPU8jDY
70VKeFfQLFL0nRw4Z8xVs4O8JY3i0SG50QQ4wszF1SVQB63up/T04nDwm4rpVmlDjwIJMvx42OR8
PcxMNlJw4vJ4hhv78rKam/6ZV4nptjkW04E5FfIedG/sr79jTFidkGvmJWkw0En5y1REscM9Bo3y
c2Ki5qQ3pODP6V4Es7nGSFcZOEeUuEYJQxfaWw5FOTvqJjmnStxV5R2ZT0jSQa5pLHideXlAkh8s
Mo6lu3MvC/tcksYXTm46sfOxC3e0IHkQMAsTnL9WyWj6tOM/CSi71RAF7DzN3fhpSIqnNh2KxJH6
Nvs3NDhhj+V1+RbMZLgYmfGlSsqP55X9xS4r35KosjEcZKTqbGcNp2XNtUJZW8cJ2wDA8f/LIzzx
iPvqBHvdr7XsERPFl6R2yQeNFcHXJLMXBqrAHYGTPbuI4bi4l+uUMOPapA/5s4tL00v+886se94h
QYXS74FSo5QjshJxA5UunzXVR+eJqlR/35EKIL8Ijz+ouCGM3h5pNg7w/hChXIIXD8MgOIBhIrC2
V46v3q5u/yLuuvbYpPCv8VVTwPl9znM3sY6BfhMrPWlB2QGy1ifXMQer7j2FDKmnZlGoSKAkPfRO
xJV+7wYb5XQxggpcK/UI68w2gsi/EYsIPtZMErj78/pPrPOgNeOZvoLBgpIQvwWbt/3yJJl8jqop
jXE7Grtk0oP6QU5TDyCpAbgUPNSypvDhfUyd2BQoq4ZSNEHwvRobgIY2b1n0gbpO8ZK/+xtW3z+m
UhlkjcNd8Ly88m0aDV2Uv5m11VDnTFXlbcPwIR/xyj+CP5F0H16wUgH2+tsbD7a1eZORHBrGpJdQ
TP51ENFPIK8/SBLKoTX9v7wC6+oBpE1TNImm6sqUKJ9zNbCd9HDNAeDxqKI1acUAIZ2hyOezyepg
oMWbWyRl6ejJoP3xyL/oCvGLEy7/cd4Y8ZAvbrgv4WYNxPwtKVvNWGSkXoch66K9eoEjDhrHkVFm
3m+0olSZYvGFn1EpIkFxJzbI+Z0v9zLAczSi9GDdYi6UbfCZUuJRKqOrKUBLuiayRzrdXqSy3c3N
18CLcMUyF2yCROfkuL8Ny85maU5dr1aMnd0oqvBgQoZYuKdMJxUut16IpMDqJXFf1pmshA5BhkAC
kUZ17fwmRHgt+qaLXPeseJFRZCkg6Xj9g9a/0ZgytWIbBd8Mg6s7D3sl8666hQzC9xoAqvs4QXYQ
Csdgd5ZDZqa0Kx+Q9e5opUtOgy2yBlVG/M2YPTLbo9ACNP3hIAG5e/cvr9Gdcq4mrw3Sw0BTJiWn
sB379g1wP3o0QI5T1Gp4bk8qerIyuWQxdHZVn0AOGH2ee55rfIyZHnaT48Vo+Ij+zT81IAv2nNRp
Opiv3DsZk+o6pLMS5ABKelUY0oCTqZrxAU/h1hyjckw/0g/qQd4PGC10jeyRL4bQfb4ryN9Xn2iV
z25jfWVsCSqz7ncNZ4igYyPKhbsRsfpRr5rJdLTDGn7uVlzNSujhmazdMHiTY1MnCtZ5ctA2QiY7
a2sxnILOdWqPSUz33WTwbfvigp/Z+vsO8nrGPdziyQvPVKuQLR7GtNp771crfNug+qkJwr9346Rg
RkI3dXvuPxUgDAcW3Zffy+by2P0Yg/7QOGPtHV5rUYPRHUGABnFlzy5Oqcg8AHjFkOP+GVNj430M
UqYbyAU2F3uuK7oKIAboLSRPwaM7xyBwAWvFZhaTbKUe2PE3JuRPQ+TswP2MQ7fFwOnnW4AkGf5e
uvZ8f4kSdj+Db4BYel1WHJl3pzbRxBRYPFSXAFOtWsueDbnvte6O7l2C5sC3S86cKcr4m0fyVING
sQNEt4tj5gGZlut0VoWGzjNFovcaedSYCkT7EJ9jt3fW7ytAV0mTv9H98wCP6jynsuW+KDyRGiI6
dQLoqGGrlowHDRJaBuUr6rFiOn5v4CanPFCJU+r5bnJMqVZ5y9/Qqp+R86QWYA4wuwMcO4GAThET
yHdGJkft84B69zz/8ClHO/uWyi+O9cNPRAkQB8YpQc7l73ASOrCAzWBVafo/JK6/PFg1CsvGkh2e
178txV3RlHUKRtkWBKcZ4GbMHSwt606RwtrlKJ/UwryWyyXFIBdMGA6QM+0LkZZgLfBEOt0gimJ7
EPBhM3YDgU03FpALzjJN4xY2RpCqJXStEoGjMfw1bXs5R1qoB742QSpS/AhXR2tlTi0mc4ykL/4p
uPL8GkpfL8UasLgNrydxNsEjoooLH7SBYo60kcOJ2cWJdzT2Oh97w7Fyl+7jKYrczcdqv3ZdneoX
ONi6Fl7xJnSYf59KmJyfMGd4/JqGW/lCI8DdhLV25dWllZxUQp95ia6wyfwix5dF/Q8QnUZMdXOm
pC6UcSPWkpt+yeKY26YwisDjwUGCtRwaico8iZcfg5idSOzSbxYbgkmUnwFVmTjl4MnraY3hHuKb
qygRZjVV/raWMkmJenuv3Fx4l9j+5/RPiT0MLSRyAy4e5a16t0ZHryChhaSStsOauuptLrHuz+6T
0XeGktSNKQxB9/hgRN9SHAaSvZRUk7pZ1F1zp/PDnoyJ6m5jsJV51BgTKZWio6ZGHo2d6IXQCgMU
McMzFqA6rOxmAqJZ0ufZTnOTNKXvUkTX9w6Pds3gc9W6LEUXNq9F5G+jUU+pk94pWfnm3QBNjWJp
w1V6e7RwoOWtaC2Vd5BhmfNSbklrk6uN1wRfMBClJi653q4xyV2qAtuTMRXyboq2XmteOO8Sw6Qg
VLgESHboACScjMJ1doUZXfbdagzIGQUnmBfIgkibURRB/Y7Mbg/PEBLSZs7/08hqvaP9VrwQLxSr
e06W6xiQWIq8ebybtcEsNcVizVc0B498iGD9nkMmL9bVL4x01+jQeh83YzuJFR3F3Fi6Lzg4lKC8
K2XJlof8zcldWnNdK2/ZCOa5E9ARNNb6Ki3uhavvZSra9Q4bndlq82U7j0i0foi5/xXt5z7BnHnE
LMhDKQq0nsN2XPBFZDmz3OJlNRs56HpOtk2t+PMZqqD8z5hxxik2YYSZ06rT/cI0z4biJAEFw1w5
SWPZot5/lC6jPKIGTtltwgsMFcMgvGo0ZVwminnt32xHoW+8nbmB8Azfzhra/gFTfzRuitwC7ZUK
46zpcrhifSu40ahcqhmRaWbfL0YIox91McqiXXk/gwdAVdm/DNDtMrimDg6IbQ4ruLUgldgoGUnX
+lmWyrEODWs6tIhPwTL3rgSCd5e4fpfpFTc1f2DF4gjEulN8P5pgJdl2mCJd4+lkRlF0UeUAEA1Y
FDtu8lI9V6RalZOadWEByzCncnnfAQRSIgUj+cZh157IdX9C7VMHeRsPEtGUxwvr7+MCO/+n+x1H
pvfveupK9PE0BwYfwSQsvws0IRwD8nDPj07y7MW94Eynf1A17e1QoSSUHVvO++hiSq6ShMuOA1cG
pbljrBWTpvPiG4jHK9aTeOTCMiLs+X2mY03LphZcctgSmHW5lgUQz4myKicPNS+8toBFD8/eVvNj
oWS9EUQMynEyrXZr8J5C9wKiRJY8KgV+tRWNCbYR01DeYke/GOJkpRjrqmjcKWJLt/c7/O7Ro+fO
m4+AdwUvpfi3M3vn0+nphnDweUG8o0z8R1CjTzClj3g0nVJR7Vi98V9gpCPNaZmji1KNjzuEHczW
3o5zW/sATu6uOE1JcDJ/pTyD2FA9IpZLBR+CBXZ4O5xO92xyAlR2CcvD1EkNBQFxtApSA8Sq6hPE
iq6YfQi06+CrHBM58XtC71fO7U7F8zIY2KPuFnSH93ozKj/dFWTX4/FJP255AuEDNFWvXkI+ZqKZ
R46IEJRXmwvpgKXhzORMbCrav95keGhHH6aZg2+LLdTL9KrHh2Ax/Yh+bqg1iKh/HmuXT0fDEIri
ZFr0bd34VEDWJfiiszmj0Upm9ayo0f8VCtg/KUirZjHYuKQzpQxB2L8wVd44L+kVmSLA7TlRSvp+
fXupZLhvxi/U9/guw7BzzrSYFE+MeBrEHfwQasO/VTvPQUYZkPi/yL9Hyh6WTRKUi+o92ugNC3vX
hHT/6sH+N5mHoICU+fDStDkcZHLmxlme+NKSDMxo5tk45xk5+aRo8+KiAN5eX+QixDctekSt0+F5
4lOyusfBRFBtvIKtk8tbx/biqxI4356grF0Pkdild4+dbAqMsLTJKig/FEaigfFs4LhQHz4W1QfA
rg5ysN0Ff+EkK5hjtU8R+aauTA2V9O9S41OrJbPr4eRZOAG44ZuixVl3MsWxE9o9KbtBLpcIjpBv
MXVESm04Duice2Rajvo0ju1QOY8kNd+ellbqLBsP2+nVoFPTc7qZ9sj321ARAJjEmLcScrzDahnh
8ZS4KOQ3svKKNMqO6CcK98U86hFW8sOhrBiB0h73exUhBHJjVBbzvgjDGUjoAxwmmsfqfqBXZh6u
d2Hx6d4InoDEutrv1x5KlLMQ/yM9rgWr00yk83mmueqChS8fJASPdC06lW5B086psZpEJmCPDrZL
a5OweXzzw/m6C6g31PvOmFHcHU0v1Jfjy3G0ou4VBwVXLgo6oC0LSSPM2D3f745EDy+tfMP03RAG
8rYxSLASxhEe+t/jc/P93B0331iXXr5skWM+u+d4eCfv+5NXZyoyOZz8TERdt9NoTfH18IDH7yT4
xGTV0dDToyR6oiFMzN1p2EhpMwlor4Pc6q/J5Kwl7zaPWu1wpxJFOBGdykbbe/sabLl/IQ+CWkh4
UKQgw0xhVTiCIP4X9Nrg4ft3VMyW8IBr0pF+b7VYjlScTXVFbljV6NBhoEcSgIIGauMenlbtymsX
UujoKnwnZVT3tku4gfU5jJuW5Hp621n2YKWvZyMMIJzas9DJzCjJAmUjd7jNcRGwzKDaV0FMVyRY
SYflHFbrTa8Fq3B6W3QVqT5R28tf5EpeEfLO7kEUdg4h7crY5oziMn7Y7MReW+7d4SNCzvYvyIF0
5a4fP4iy4deGnqlDmvwmgy8BZW5Db/CMd4ggwpx1vu/odAqFi3P/2CphWOS0jUv0l6hAT88YVmzx
KzRtcV9HFNJO4daFSIe4hKbGxDWWkLhnugSBYBBTjTfrgFGBNeYeAd+P2kV8+ghCRKCRvO+XOXWg
8t/XiLz8MzJuhlU9s2Xwm7vci5jzJZtP2a+MZmtcbyJZgUTg2HB8RfZreR3FkhJDvIVCCPyoGdo7
KeiPtZgpy+MEWEl1o2s5Ii80OneQZakhZJ8TnHKoBNx1akCw8Z2fV/c8w7u6SlKDfGehw8cXfIUF
ghkihmFG1Xgbs8SxN/PwUakhsGG0EtsT9dLiqQR+TBJzjJWux4noFk0RwChYKv87s55DOVxGYPiA
sAejJwEM4r4lEaRkCtc5bjUSQZJb7BiHblG4dUdAXilNMxqrzAkp57wbC6+44e/xNoYEoUPEHl/D
87eQXZuHmog8MX+QmSp0+bt7H0WSTiPgI0e316C9p46+4gUNuI49YS83ewQ6X5sq8dbiqar5z2MK
/I1RVPU/Og2mMcX6Cuy8ySYs5KegyVvHERoReqTI18+bg97BdAKfzmNTqIgKY9IFGL2Z1RsbWDL2
AFQok8F8VYoyp3UsNdVvph0z4KAmW7HV2pZIhzK2qfvY+273qGWAAUH3W7c5IZFr5izV68XsEd6O
K8nggg84eKUBlGCCenEp+aB5gcp59BVAIIfJEJCT+bPfyghkPAkP9VXKvCJPwVAom3Bcq+SO1bEN
oyHSo4lsjVEBQ5WiEBQ8eeKuu4I/GvsXMa5TdWDlK9c5ZIZa2uvQO8DWg/q2ns6gtEReYFON3jj7
PXIAH4TYRhED/J126bUUwOwvUMCjj80Rl9WMgyR+I8YaEf2SN3ddJhKdoxUj3OWUHjxYIRMFzaLn
gifrOkrvCP2lJheq1HTRMacmaW+pKioHnt9Pc74NVeISEHCbW5HFqqpEJa/18DZjWEdE/jq/XN7Y
rPjrs3VuDc6MaT3dK05Xc26fZkV7Vk5qpf/XBz9Unmp3EpkgVDGt+/cVCdIbY4gAIpMkHox5cnSM
CQ9OAbZspVl7OwrKYCLWR/3F+pS7tFZTAJN1ci1EDolEdq8cjelQygy96i6O+lXEnLH/mkAlv5X1
AcR1T1H80GCqF+8uryLe2CuunMnjUVO8ygecOayBqeerpUGbTLdMrlR99eYNgtVQYBgxZWsktPAa
ZuwJZ9SRe2pVRmitpZseZ61HVW3l6EDd13jxsMs38C9eu8XVAKaj9W/6qJPImG/QzWns+DOxZ7XZ
iT0/3VZxiIgikihcrAv8JTLizoTcKjkRSuwmligyNJqB0kP/L2UyA5B6IS8mWC+E8GwbkUIOuZ8z
4oMqwLBm7e6IMgfu0Pxd7C27pnLG1qMtMJYxOiFw3u7PNpm/qqdtYvjyEkD625UwQ1KQGTTCH9My
iJuMiv1uKFL8uNWHlkzYPl0kNL7a7fuRZuh+54YglHS8LzIUoHphntd0DztRfykcsCPehenYi04u
0kHFnZ1LAgu3VAnFIBbQGThPVKvxn+hjdS6lZg11otLpjeJ2kWN74E7xPxuQffsMAMLEWdW41/y5
MWm9hoQ8bc1c8RdYT8ORSAeK/u8Ga5S5X5emAU7LIaKelaCX6f5AHHDyabee+/NuaQNaoP6BiAMm
URxnyNJzgziqGDcpSGyDoT1qqy801xGSJCBB3lo1hN2Bxhv1lSfmhY+FLShS97e9AoZPysxCVkJo
LN3PHiDkPHOVPc+viQp+T5BEVioWlol1rmc3UCy0zBFPnBySE2DTnEoez4kOrYZSweXdLEdcgAep
wR8+utDFvcubkJ9B7r9prhrbTXqWEJlBp85fkKFlFC9aV6S9qnbRZ3Yho4EWLiUjEHufqoZ79xag
MK1wTs08JVKuBdTMchJMiQG8lfHcc0qp3WXVXRSQ0JSZBl+uU2IqljNu2tzAIWnuLCooj8Xr5vQs
J2gIgymTFM7dsj/Y8OYcXLi92pzVCasH4XAp7kpLkjl5xydSw3LY0tOZfkyjlgd91TfHZslxevNa
mnMY/0cwArvTRmghDCz7tXXh5TfIYo4qW4tMI9hhIOtsTjVHuDm7sw7x/kwuXqUypRcqDCNyvwAd
52v9/+rIsop0L3X9Uu9CSlTjR2/VKi6qgDvXVxqHLMfstly0qCYKGZeGrRGXwALLrX93y4NMxymY
7q0vfJ94ZIL4b+JGM93xyVh56UY9KZlHW/cPya8yUw/xZYKMHEi7i8ea+S38I1R3dK6rBk6sbx9o
GTtoSA55lu0ZSJVITXRg6NeZpomLp6K9v10GaBycyvMFrdv1W8DtiGuxGW82fzBrwEGw317ty/uz
9cJImmaP1kbcDnLS+OgoWPLeJmDNigRRj6V4KLT1oDL1N0CqKtC6UbFMNeuo8yR0dZ3e4UeipxHC
RV83BvVh6VGckf56Pw+ksMNozm6wvb3ui97NxjEsgwYnAWjxF/Af7H8ImspuP2JKvoA/jZVZKCPy
PTFKjYi7mcSo5OsEs/avAIH2JqG/RVUvjvn5JDY5/B5ar0oRKjyQBk0Qboxv6PAyG7eT2eqvOC1H
Fv5V39SsOmHP6GK9FMI7cAmg5fEzRCUj84l7/47ois8uuP1b00a7HqxUL0dyYJgHv7y8ye5pykl6
6aGpNYdThG8+04WWzcDnc4/4JDPYkQw8Zkm7gKpK03Fscp/26WE/A+sEn0SidWwDm7Vn566ORw/+
AJ/m9lrToTPC8EnjjdwhHk5TFPTXkZ6AEji3u2kIvhS+RZgMk6Ifcd3j5VupTKFZ++Flej6jfFyq
iN3yfNgsUBj8JlGit5FcFve3dlAaNdAwJkWasBqcr8YdiXZP89vycfCQ6moru3FXlWuOa+D0w03q
jswdghMSZ4ceFIzCku7hx/t6FLRCHkkIlls7MohTY0k3iQTEsDB/hT+Fz9EnF57rrmeKj7EqjxHS
Ya2VmWjlLFIR06atRYS+rhb3QX/KZ33ezNdgCZOhnN+UwCNqRnm5qFS1zrGGfLopivGSzX5TFuac
1KdogglB+VU3zs98fmmrkRrxWqQoeYf2BsQfjXtWi7T0UHdO2THmc7d7IfBPlUG2UzOXJaQI5FJX
5tYWrOhXfISRBpVlftXUJl1dO+e4zF0kGaL+TxFdtUb22gyUj4R1gFRFuV8DxFVMrHXTGARby2OV
szDX3oT5vHj3qi6c3RILdXDh+KydpTCkzyoqkM+kFMkGppeoI5wPVt3Y38Mar2NDgSKQnNGKvM7Z
Jeb7DzROx8exBaj/KVFKdTvq/XusDy5D2atgRroUBFNbIF+1sSPxxLFkv6siBYXVj0oYgYXYeBz6
ObXPZ9jvD4S/RXOnJGPU2mtvKlkWQLGGYkNdwc/t5ebxZiWzo0deis3BUANyHJ5XD4PmBlK/7TZN
ZAMifJP/txVWIQvDThNv4eurw3vdVmTOx1P34OypQlrQnKeuwurgUevEKpEntcAWKO8vbAw7Vq4f
0n7gPQuEvybfu10I1EoenjurmJFnqlRu2Hs4WgA5MyfMph4C6vqv3AYC9TBO+aJ4X6kbl5u0Q+QW
9WbJC80cWT4TndTqx+UFRPdaWF+Paoq9xtFk43nhsosuRkn+KPHMQnBOvu7+uwolAvyj8l/qgxiK
MQigAyzc9ij3m7LyryaZHIm9Shx5Mcao4QC192aMLx+AwtrP4unTGG1uozJShErFK7wpLxv+Twtv
CjLT6xEzKnI9dswsyP7jfmtTchguXNFj/uNd76dwAHBgZ5QPeMWhELH7L4HXMaTiffNH8wBFhOMM
DqCUnRjMII+St3TVFPCxMgiJA9MAovRLqcO/ivX1ZRvcGDPwceJDTs9C6YxtA4gZGW+er/ZyquS6
+F2kLxdDY3KW0HKF/XuQlAuJ6LCnt1nDFRDUXJEnOSzgfUmXrKpRVme54fQY9cuKN5sGZuk1+N3D
F1600ziGWYvCeT0/pu/kKUDFv0vrf7YNlQe7HuWy/H0yNPNPLyxVp3v+89zcfwR4q0F5gaSciPPr
DjqcaEWVRfAdSVil4x70AHs9Sdy12jt3pmDnaM4BwHKECkjxD386nziiK3OByD/A+SKIYBgHwUAI
f6HHbmXCg4G63sDXf0LDeR+jF4Nw6Z4o+CK3vuewNz0sp5b1b5Zlr1yeNn1XWa8rFwmFI0+IjmOp
WL7AO6EdK5+paB36U0EXah7OXhmrhafwJo4J62Mck5jXPzd1k4UJJEqgZxqds6peFr1czemsaakA
9GouYO/rYfBM3LElzjNvuSRec8hhyWVS9cSR/MAzUUMkAmkODNkLcRFiXQu8HXTbqS8EwSr6luM4
p7JTDmHvlBR8dAeqpUIt0NjRjLAc8udViY7KnmBo3Ve557uNShB+1B/4tZEaT072SJ3hHsiaCvlq
PH2chk11lcyCwUPPdYG6K9xY1lejyrxDHxBByXThyupHLg70Eq3Pqqn/s04VzhuF6rSwadVK5m9W
SZXxdYtr6nDoQri1thLFpHMPjJ4ySNdk0dN8KaQ99CCN5AQ4ttzEGQrEHYHvO/twCsMX95HWsCq7
BY9g102rMWHA3mOKUSTn9Iw6whZ1x60HiRufQ4yWD5Ne4HASJfSsAyuhHtHoDIHg0iIaXtEy+ZTs
GT7yWpbyI0dZbEO8khkYRCdB7IL/8LKqFygulobUr2Hx3e3738B52okScdKpLQxqc+tvC/z7GGfD
Oyr8yI614wxj0pjFzHdOZe2HopZ2hiFKcBD46Tl/A21U+IDeOvKpyPh6y9/SrNzLvzNzbybAwJIH
Z3F8k+vzot6VXvNidIt70Vu3mAujsUgXL2b0um9zsw72XkdrfUWnc++IffkvENO0fam3rHyuTqIz
rwsihyk0l4uPgPEaGxqDozph14iM+3TZxV+whc6P+qtuWxFGFCgfiqe4fLeFRBOAUDwBmutYGAY5
lG50VBKStqsjPBWTD9vHn6M1Otc8K/y+I5ywtjUpY45iK+PaudIaqTNJ31IiWONRXdK1f+86hjrE
tkmvxnVYZ5jkG8gIaCReDpAVSNXKs2wGF03PCuBwMN05lFWwDZQ/7h0DIMsB9h6olVcp3IL5FgCy
UvP1d+1wpgJCd6ah0ESwvQ0LrgRGNi4UHeRdZ8kB7g1uP918UaVtr26Y4MRxCnuzHp1WOKkQ3yD0
fdOxsPjDdRXYUI/yNNo/8ERrlkrgrOdjnLfeQMnZEb9dXbLH5gS5N5ekbIei6Ma/IM09qZJawhUD
Jjbe7axC2o9tudmC/TdvtOjxUYc7wg4016sURSryPbX/xdOcSinYEkIzDAmqrkLXuJr6iw2UO9/J
1B54E5c7eopUGSRIni4mbp7juHR3K01sEtY6NQh2yuUS6UPPvRxdK9t3QLlUYNIRNzMQrLXGay3f
As1IWluiAKvmelWp8rjNlUldJqyjrVwlcGtHk/bqzgFOgAUZ4MT8etqnnyTdNYY1uNP3GeGfgx99
gdMFU4QZ4XirKt2YLdlvazLuvytHAKwS5X8MSGh4pzDy8wAMFCI3hZCOnbJIMb7VUP8Lq4XvDzEY
N6jxl/qW0lbd9pf4lQ0BU7by21y5K0DzF+dT91p1vX7YXWRVIpvtT36AlJjh0L1xpWHMQcHUQhoz
blj255cTS1P7OrS/+Z72JDoIvO7HcCRlfzY2LZvbr92AyKF30N+s8RLqfvmR25UyErLIN51KxRJQ
8+sLw7JaVnQRwNOlJw/TEjcXq8njwQBaRm9C0agHMeIqc+UxVjIFYvBvTvriezhbQDqXuwZ6V2e2
ilZryBDjc6TM4wruS+qao/xzzIBSfeJa+828MYmzYNvQIf0sWwCEDsW63MWmuj6XJ1oc6o5ITdcn
2ql0OWdWG4uGGao/9H6L2UE92t6mA5jN2bxiQoq8aD9AavLci9IcUw7oK8N/cD+3ru2MvMDaNyQS
kFXRFBwF5OCMl+4WGiRuHOUbXnrnDGyc6LLadNMnrsYQQnxXvqXR58aOUFO9KXp4dwTu0/2n1ye/
G/23yz7EhvH00fbsACosDCjJazgQpjfDwZbiChwFNVKrPnPQzZaS53b29e1TS53jGfFsiTV76hy0
wpl5lJj7HUPMOnJuNGVoelaOc1EnykCsgs1O7mnYp0OeeTHSm91WMBrooZgxsjxfSg855T0ojdnx
N5WMg1+UtvSvMAolNkSdQcTW8WaJrYvF9/kPfevfhSHa2zk2P5TixB0U479zKAz7GPOhYZy5agcI
y6BoXvnnDTiTq7zp0sLlOyyaCk1x5xz3QpyF4EoiaKmY+Hm9fE2bJnmjm5Do8FL0F5X52gOscaF3
672TNejoIC+JyVGKp40U5Q2J/AF0Rmfq2vGpgw8PBZP0At1yS+6iyuPCNYMCVT9mdvX2y1Q0NVl0
em+la0oPwVEnYpd9joBzJFyYUJTWY22+yGXfpX9kNiZrrvEeICBFTWgZKV4Q4hhBvkzrSzxvt6QY
MB5A5uz1eHFHlnSaScu6AI6fW4WfT1kCPm4buaoIHeEkzoT0uIj9LugP/O6t71Xj1DycFWKYkIca
ssnRQGVhlPxJpU6PW1AAIj1aIbQJWdcRFlOaw1AGUiNbxDp8Iu80vVEiYYLc46Xs1IcntuLV+58z
X4pUglzbRX9RMU0s08w4gL+kp+Zm4AIARYrGJKYEjSo6U4YibAkvZXD9NNZrjmhTlZVJPVjgCT5S
KEXPhixEAiiv5nFhHSECHTinugdKLcX5a4pIy/ywhXcbag2Wo4s/Hth9uW1df7thAOmKj/rCcIf/
oLZJs0ZVFrElYyb0+XjxJcXCXmH27vyTwr1h/wSPVP9Ou7GFUvkVpwRQQBDwjvwMo2650RqfU6ba
RWNwVbm2qvHOBQpXJMZMG3MyYY43vHBxCYq/Nf2GeddAnAAcytmz/OdqLJ+ouuqem26CU7mIsCHL
hSVi/vk1AYVTep77mRyGdgIgRx7fxrWndePkb+USTc0HeeOw9ZXxmlNY9oK/nb8w0j0tsyQ/R4+n
iozQlM4oBSptTepE6yIWd7UVMaVPFiymLSUin0+TF1d78ehtUonQ1TwVN5hR0gT+IKKqvh4yTe1Q
iKR3Kc6S6+7gOn0PtITnFkdZttRNvPcgfApYzc/hjGM5d+5NSWnkU1enoCcITidO26xpzyreRapJ
CybY8bBOTb4pkmlPrxZM9dJehmBtXH9anN0xcigc36l1tTz6Dsao3fTR42+EQ+DHCR75NeQ3JKkf
JYHgxHDgxBhk0G4XCP+dowQvDQvd9WZZ5GkduhhVIsIzPhF2YKAs4S4xvI0U48iWHPauO7ppe+iX
QPqt9oSrTjyeufpSw4VFrk/wVTkHYPl/OYgacfANdkdeeOe3fDv64SqToPUIVgR2MjlKYYvZq8/E
NrBkHsYjGon1X2+s9ecEQvSFxtCOs29l4u7arkY6WMo1olrQmeoHlw/P729DAewr51Gi4nuwjh+7
bDDq6aVOrm6ludXEFGajutH0ypuC/groUvrcg1E37gmpTsmG0dEY9EhhXHZGQok9y8QQKsOROhbz
TtxTUd/STvMA8mv4C/O4EH1g2lvWMfi0mXl0vMK14zX5D6eNSdj8Tq3Ajo5+QPqjuekYZphNfFbl
LvMuScMUghxRE4wNTSkNWWku9eXkbhOqMSCic2lJQ3PYtNexlExtH3gixZuTrH5u/Y/gv2Wy4TEq
5H9287W59HZUhYM4PdfqVo5xXGPv1u+sVd+RftvM6d3RdEut02O3gEJpYuHZUOKti/nA6imgM1Ti
ekL4mBS2v2ZU3Twtr0vPQcmWP0tbXH/tnDDjgjhJK5NF/MliQgpEtrwuCRkwGX1WLZMUwlR2HtWs
uG0Otf1G24yjESBCG7Y3z+Oe5NJRb7j9bAUn28IlWDk09gakjGj2tUL8MbdesaHPFSf7Eu8EFfWY
JtbNjSaSrY4ABHKlEuJfDCbvGlCVfv9I7pFWYmvmdJ9wnRCO20a1q9fxExByxeuRdbArjeFHYZJb
BfuFpar77d0VpnZJiKsYbJ2rQs0OjUmaSQY4+1AamxQvYZ+G8HsOq9GKJLNxhLtwu8of80ca6w/h
7fhcD6S7wNdtLsL572sNh2iTFTz7/r9LMpyNKxgaRn8Lgq7TuWXmYR4oWM68MdINbAlSW5Ug51tA
r3BWLrclZJ6w37DKelJHXNn+g6fg9f78TIC+FA5uVpmVkW36YeNaN1sWdOAVMQLwdtSY80YAEYRL
bSjgNw1g7K+QEDdVzBEoFgqGnr831HmHhTK06DoLm8PeMmKmvKJXAK98L4D6rbAzhhpLxzPtANYi
ZtbAlpxvz430yPKLJWxfi5GW9QpjE4tftcou7vauY+cnSAJn1HBicu4+wwOgmYrprZVY8U2VKolP
9xUbTSNWlN3QbImeSnILKWmYTV6YiBag7gVgmEcn0OxOjHVqXH4dOfudeszBDfYDGBGKRT0emrW8
41QNgymDmkChhv+J+kpO2qFjhQ5Y3490dYxwPIv5TmtnIce9HWAzbWVYNLHXBzeggR2lmZczbBEk
Z6EgG+pYEvhw3/6qQ1CQflEpiLFVrWbbNldnygdrdraUTXUcw9+yZGwEcdQN4zqx6fSijZkXsWxl
zYWyz4B10x1Y2/UmpUmCnAu57G5cEk6fIhKxdEqFUDtfrtCET7+qyWZS6uCA8jYwFG+nvyLb7qmc
vF9iiGI4o4sFapyaqo2jYS/JbYgPMgKL+SAgXSXyofV1HQOcqawD57BO5OiqLzdR+3V1qhE+w2he
LqEHrdzAMaJe7LfOhvjFoZzvr4FPmkX/O0ty12Ie9BaloDRm5r88LCYuM5IH0j5cr35747ZIzbkr
+CeLwZ82aHlnXDTprxaYp4k11ra04Sx+y90eU490UP5TX+UrdGuzrCVnT1Sm+cEBNGATwdvYiHAi
KtmbwuesxG8QGp6OhkcnJSqvbsKe/c2dGbr6Sh8WOWcZYsVL8cT7fyXddKi7hT5gH+U+b/pN1Xyo
Sx/prOnPWh9sFkHx6bjP8xck0rh44fW/UNfVC6dhRy7nC2Mm+JIzI9GN62RxqQ0SRHh4/q3hyhNh
Ic0Gt6tF+CAKE7jRbVLaINzlSvds5pqXIZjUtQmI6UQ9TvyS7e7Sj8/uAAnIdWbHjMm8SbULSQTd
YJVRFwNGUhuwc/Iil4zqIpUgVzzFpwO/hyeVghVT6PyByw5oaDqdQLbQfyy6OKGzdNGXuV17ftYE
SVQpW16GEXQ3VtHTgbguOdbz1C7G4rsVnlWlveDuY77GXfi1NcF7Begj1R3479QIXIErVZdBW5A8
TJvRzfvrZunTIvmgXt5Juw2dl1hfXqxXdC3M0l3K0SODADaVEyt5tWiggp8ea+OYY2iZKOZ4qsOE
Sjyp6D7CRmEbmiD0GOox6v+D+pXEdK01zwAH/6AumvuiZz8tbfK+yh/uTEgu/Y4TR6p0BDr48Vnk
FeK0IrqqzFi5akbRwFa5/OqnSEXRF+svjF1iDJUeO5YATrN6TXa1DM9tKDMBj5Ov8VmfSKxUwxXk
1I7+DQ8age0MXSSBkanXAA2Nh9mXDrFntWsBQRym+a+VbRYdrzkSboomqV46aZJlVsqRpfCcXTOh
vueNtULgWj60smH/zZY1NY6Fl+a1C/WCOX1PG8JcIyq2Oz1TLZ+ycCBIokYj7omzdx3rxsp720jB
LFZSsVfs1iajbq92XYuDvncif7ydRtPeQAx/eAaalMvGgRMcezg6NsXMbmf8EOA0o643YBXkY/jl
4axMUgqfx6ru8GD/F6gTosUaIMq2Eo/OaoRXPJSlu4rYTketfnnnMAbq/J2bWH49+vs10BRc4CuC
/+fhQk9YxH9CehLkpBVH6/ed7WmL1OkW58m3ocr7PK92xQVfo6Bz6Ti/rO2vFOWs96+IhXc4rVRr
e3H29RjrQDRx7yMD6orGxQsyJ86I4r8OiimltrlrLFHpoDavSkQ8ae+ijuloWbamoxoQA4hmi0gf
f04Cx2iWb44U3nBbDLgb50WAVPNjk0bfjNIu/ApV0j8aXSKJTV3U+OVNHG+RYS7oT8AY64fQf86y
07ScUnhUQcY0/QWr+gQdNU9Ivstaj4rmhsHSyI+hc8sehWqnbocreSBtfco0EseWee5CH2rsC3Kp
91VZI6AFTFwVGtavuvAsC7E5BPBhRXi25iqVI1dmNjsoZSXbn9b/nm0xgM9oyu34o3UWGZU3bN2u
CYoDgF9pE3V+oh+/QXfv3D3nq6A1NHNi5iwNeHNqtdfg37WNuYEJneV2dZCalpLZKHuehlGTmly1
2kta7SR3nLASGbhDGnG0vAkwf9m+kTl1R0DYWBEwMw7zRJFKH4LIZA/EaOkL2Jez2mP1GK+x6XdD
9awAk1L28MT2ujPsvj4CO6n4PAJ7eBXZbfRIIWcTvufkQoAWZ8cqryyg8WkPmBfiYUxs/fHbgRsq
rsiH4gQtK9xd3ghvYyg1J7jR2BEsFofsxsp++HxIhMj2gTjG3BitY/hVFD0tmGaDOkJX1++uvA4k
al8KZ/S41V9dctiebY1+3njKPDJfJTcH66OVs3WicXj4DqQw3f0TtuIYKmicvivsFKk+NPJ4Pm4T
Rew+SsSVqvnzCyHxR9I9B+E4DphqVX+PG+GwMXGMqC6myNbOkf4TGaKrmMCD9af7wWZL4ZamlTN1
h/zqrgO8JbRo6ZbHLawCSGb3I8wCzko8lupm7w2+QOX+dnFl1qjVQpTMd3mMbahtT1mQVmgtHSOz
FW3yhfT983Ab0G+jg/2iQnC6VgJZExPiheK87sMp5gnli3B5Xo7iVtcD2ztY7Ok6dJ/OzKAMprUJ
vk6B1Kg5/bUBs3/mWf79Qcqg7usnSauGIVEp1MHazISw52iHJ+JMjjsfE01UDkm2WfgkvyOYJVuD
7ag7yliBR0AzQIBP1KJ2uJzvUsBnieKSDEo6H3fwTHz+rV8wvGK/y2Op/+sxZNQtM9i9X45hMPy8
DAViUB4/lSsO80mYPxkE3V8sOzR2iI9EUTbGOaSHaEoBLNWnm3Xx9pPwkfYrUe8CA4LY2DuY9fkr
olqERcPc2pJgQJVzl9FujD+lRjQoYVWTW8nmvYLL0XvfuFgAhFtc5o+iB39atFClROlRrGcJmvg+
/a3PKiigHAezuq5/QEWIS9tpAu3iBw/vjRFCbNPUSrStGjfLGzffDwOXF58Qd8QkPyTYVfpogK7t
nqjTPWQmBIEM9s6kaPriZipdbDU5YzI69MWt4NLR5N10UJIhwfDypW7+qTSfseeGd3f61cZhQW9z
/p2oCkDgVw6eE73Xbqw5fn/9A5KfrZ8WGzRfJMA7wXkqZqx720yf3aAZZ/CJqDy3yl5vZVjFdpj2
rOA/h2M1ApVGCU0waDjpAtL6uqSsJORDBjuedr8oZfDnB0vIb4OvPUI6y0uHiKom0Brx774DefH3
RxBVGhRSabPXNn7/mTQUv8V0ogEEou8ZevEmy5rQNLtV/LOX9nCCxbjyALLRTUs9JTulqq/T1BfC
GLSMUHAyASsQcltBiB6bS5bpX5Cw9A51y+R0E0EptnEX4rzoqFS6NB58oAYsvBLzzeZCM6SZCpA1
Wjx8aaCwOe+4hlYCJ3NCrUUsv1K/9eY5QdLEADKP+ygpzb7WmgDytA3LLmxri06mCoMDIvCmo3rO
l8Wf6X+qQpIs0kWbOjy/yfhmPqIJLGPZp7EZXtTURvpoHa8mV7cPOiIAirF+p/odMnYHB0eO/b9d
XILnqoE/egB8m2u1EgOL2mHLuIPr0A/yRp20uhlrnqOImVMXGh67PsjCXXQzSNpw3XSX6/AcZyrT
kNrFHkpkS7gMRuA/bHdIVU6U6JICB+yq8A0p6kRPK48SXSNjiWybHx6Za0k8llqTworJ3t3EOceY
/6ODXJK+zFkJ7WBJCzbkBbYEWdnAnf112ENmgxLzVjY0UzCbGjdwOeSFO/a6J3Rxu2mzovDKgPzG
M4QCb8dIm4HJE1FeDATX+yjbf07wGbrdU50gzwH5irs7W+M4sma3tpxJtL6jkNHxLdiajQzikpcg
plDDFXjFQPSYV/QcGZmcAnljTQGF6NTXuG8C3jTUkL/HEen6H2ptBoBzPjCuiwP/7+0d45dC6xyT
bzFv/HlEe16C5pBOcRiwXpHPO0qPqs6dMmuR8VY3UzkIj1++drU8d3xdXPYM+UOJvtVgL2L95z/W
so6sbyslSOsY+zDE010wt3pyBZRoLZJchFTXcHkylyoRQBIayanXafguIoUCMtb4cgYNXwGFebho
nsEpfuWkHtHZuv2HPfiP6bwR+pkgN5E+OZL91+U2pw1CvILrHwkan2Zzmrob8wXPilr63ouZR1zk
0I5jeuJssiH0+VEQCaHVHew9bfrrO8iqo76hd7k4h1yxX47/ahrlxvxY0aI3vr3QBtY71BxWi1Y9
4Fj5yI6byZ7e4sA/ZWCbdxpiBDc+5xN/KijsDu1h+fwGmd/NFn0D/FA6jkRzp8krCf1EZDDFMPnt
tDXXK9XprWmIwh50zrkbrVmASB1TQOdzu0BBdm4j/Qzx8Wsr2287RSXrwCo3u37o+Y88vBGaSZqL
O+PKHt6m/UwZkZiciQEx6nBqzQR8N/uHyGHmz6vewxJW/DmHvTNaVEgirvCOwdDr38L6caWjHFti
+ITKosDPM9JnMRIOBhQN+hBlWP1LYvNYN2ydMq3CKk9/thh9ysOx1PZv7wof3Bdz6ETG5Hq3Z2C6
x5PjXdboful+VyCeQQiOIYLSfRTranhFlRgLVT3USYfQXt6jwSrGUXnGePy1LZVyEJu6MPi5UYQi
2x1F05YJWIiWyJnGGmugvUKX78Isl5Fe6Mwn/OXmPZmRD99LyzdBucocUFFBYTZR+Kt3EPXfLeu1
EavGEP0vZwjFsXNczzSpxrzT31zvLBpBl4uSX2zyoAT1IwLyEVmKEqON60SpCxZkTD3KYXEWf0mk
mEAfEkJTJkjKtIsw03cLCR6B1zacGK7hjpCL+5YCBLxNxfm2Xs7BI4h160idbkeYomEy5JWESvTX
RASlOiyXPhrVmlL/KbI+7Fw2CCzY+kgk4lQt160Xw66Mi2cVXVNb0NDK4lQSOiF9jYlwm2YA2oFp
ILlOSUDtPEJZ11DbQmXiNVO/VzrPgAexrxIXmWpg4cfDhYcNNjkigZoR6f8FtJ2taatPgDVYni4P
NAnYtKf+kaaNOw/8c9kys3oDdRlNOD2aiI7jFl05SKEenEqaZwMIVN21+zGHk2ga6nBHe0+OmF45
10nNeejbalNeX7BXQ8UzIXR6plgKxFgeEsN5JAqJZCKNhSYswz1JlQrPBeWOuIb5k42R0dra6T+z
hvEBg9wEumW3OymvxqH4VdViXni1Zip/8EZJvueopPG3hRTbGUZNOA91Jr6ejuZabQ4GTMIMtS/h
TQpwaT0FMsI3W9wr3BTZFDWvEZ8fIsfzm40pkjZFbsUvYFX6KO1qpSUbo6S9onHqCE0Rjm2s0ST1
YEk9BaWhsoq1Oa3gadbYnvtMY8OA+j5suV15aDBrNc+0EoFw80mm1smGwLs22dHqlMLPHU36L6x6
P6k+kxVbBuBPyvAfjuuB+b5X6kDr6vPKKKhl22BdY9u0CJHbXWXZ+kqomJJUGVxXXZ7EMNNNhJEa
0yOfXX9P2knzNEa/d0kGWfACjlNno8ZVbcu8cO4CzjEN7F1MAX0HAEwhScaUUa/7u2fO+2EDUAkv
vF7gIsa2lJbqukqO8mfHV7wcBHplX65eVEChyaC19lwGBdIc+SKby1D+sfrENmiJusjrd5nyw5U5
cA/bsOj7EAS3h2pZwwIiNDtDQ7bTBYobwjuLMDs6b+wKrrt7nGHIN+/rjit4SOSngSUIB/ydTVcM
/FoG0m2mUBpJZhHYdcah3+Z1wmv44QPA5ohUumwaWz1AJxSmk8ix67X0vDctuqzsBz4FM5/6OCxH
ftZDsKLfTLmrw6ArhxfznC3CIwkXw/bvXin2Uxxo0hBAh6w7sGQEOwHhS2F7+9K97TVQ/SwRN3Gb
sYkT8f03sBbnPuPdrQnviEGZjT70vCg2GpWL/y4TW7yCKVHf3C7v7Zy/NK4hzL0F2oz7veKkUp9U
KIF3Wuh9DO+W5wpjWVX7/AC2DsEMF0ymo+29wkl6t8rtDM4BsYkjcYQZZWUBfL5kSewK77GKavFf
2i3pt9sqrLVMlnDpkWYdUB935UB5sEBLrlp0OmwMRpXAVW1Z9zFngiTGIhZrxSJJrqIjiqkc7WSZ
6iaKK8c9Qe2DbL5a4W6ZGMK782R5ekVDXmOYrmlNjAz+DOhKqC5fByi2B952Q8sbjhvaVvebnIV2
BL7loQZs7HFZeW41W1ounViQLYypIyqkP3JlQVuRSVCy0xbngS3L1AjjUIRLxhxWMK2xQerHOURE
z2Xl+Xxv6Dhn2f9vNWTGkXerYiQDEHw1TZhhGk5tA5ev0d2vMFPsHyge4PK2LiEOFoC5eG7QJgH6
HNA8+LKv4mwZwu+ToTmrmsRgw1csNc8o4ZI4RaBd4ZDDMjhhJOHCNTQZ4+uPjXem0hEMYXPxOsxJ
NS4PZmyGwVlVw3yXvimY0Xz4bJJPx2OJSRLobczJtc9dB6VeGPofXsj0FFAPCUFX1C9Av69JzqFW
Ne3AMvkqHITuijUcGmi3cewUh7D67Uqwq4Em28AC+DvPmYwHFRFtWrj5WaO3fMXEi4YyzIu12qz1
CPDsKH4r6sMDF6QpwewRMijUgehG9z35XdXkw3YlTxMzfAyjK1oiZ6YBHfM+s11Sq9XGg8P1jUES
oTmPF1WaeJqkdMohjbR+89pnZhxFt0ABQ2Nt4i0XSo2DDjFJ/O8BeSQnKPQokDHlhrBGk2vOqBuN
GrIb8VbDcFSqZxjzJ3GKQLenMHzpVJEvL20AXatbEIw2GSBL3KYNvc/2ZIX2Qf3OoapywGagr/N5
kpwzbssAsXj2yKlPqaZNY8x4RGJPSmZUsC1Mc2TvL43jUdBG4yifKF5J6A/qckjKLK6Uvkoos+EY
G2LDiff7B42fPp2s092fmm0zhaQkfV4eyn6aDXVBBe/zJtRpj1BEZJLl12wYCmEuR0Nm8IR8cjah
t+TMmXQ6FOubTKt79kKYknxkvH7ptORZefsCnovOT6w5MNDvXIFM0/TGVcsGu9Cn8QkgF77VrLo+
kFKaZtH4zuNbjFL0jKGyy//rTz5VQTQoZWTe1Zae98cyuwV2jRZQrDuhbVMPRxjBQwGAvGmh/oV5
jBFpToM/o+Uf7BKpAIiiIcqKsToj0hoEkypgoLMvDy9yTwdpk5HR2iPyKHDCja+f4RuBAZpJgu6G
8plU5cGBwhRixEDvKm7dUVlyNm8HB92sSn77Uf5EdwQ6sry35cyvSbBkPfbz3EQCUokoxG+pThhE
3+GhT5x4BnRTZucP/eBN/7CjUr/Sh1VmJuKlAJ3vw26rPhfrsMtCIlEjUjwnEokNmFHGdUbpwWL4
U1Os57rxiA+bYiBQofuZBdIMLqip+prsLPqYCZHUpsqbd4MGc4v+O8n0bjpv75WfO1a5yMdBMV1k
KqLhfQiwC/FbcfFYqod0Zpf336B69Nkdhv44SO0wrQR+jmHOJU9Rm2SMMO0nSLoH7SWcLtB1TmWA
jqhGV3fSIzll7GDmlRuqVKxq1pFKN8o6eJuUCAmCR6qHMB2wSlhkF+/wZpmX/7CmvhEUBFOg4kHB
l59Aqa4RYSdeBep6uNTkn2lzn6Bxk7lXFRR91gsYFZEgpaextO1wtlmeNLgFHesDfqtuf/nj5xlf
pQbMUrzSEQgcnz7+8Rc2m3CC3JQAS8bH3n/Kb5IjS+8nwbmCCngsMx2pW6ENxCbmY/jE+EV72jLg
oUghMRgR1of5OE0sczUdOAhPaXNYLMvlefpA/YC1ZsrxZr4dBU7GeTACscuRKWgpB3b2C8CYNPJq
09GHaAmwt+8Bow1+pM1R2RI6zZGdXIXoCuKP9HlLzBgUCYcUWVZaposzkBH7DaWe+XNKw0LbDXRZ
Wr5/oQnMN3HwwFxxCuXBbg3PdoNMnr0GiO+2xjegPZn1AmYS6YfTjPA0xM/7uZPzJmFoYnueXXTR
1/I3InflmjtdyqMyxADADTL30WsmoHaq9qy1yQ8qXHK/VJvobBuxA2eHJRweWn3yxud8khvBE808
HfaC2p1fhEN3IqaGOeyHhSJMTtXdxZaMABom6dkUaxMcDxK6HTJzIEduKi+iYGLwbLzyJNnlOZ1P
eLTZnb1xY31mofrCpAUJcrQh9c04GN7FRFxSdu4HP12h8JJUgSj6iZteo6sbLwJtunePdvpbpVlS
gSM6/2tx8RRVRnNTOkh7WBF+NgXAJ3mXiDxJl6ttL1hH23zr0IMc7Ak5LLI20DVX1M8Yu3z+aCHL
MeHlwEZEu4tnH3sDHMC8B0hHRnJTL8IspEwFaKZ+PP6AIlLqHcVbzTPoZV3mKMVli5BPWhtPtWSH
0SiZwR+E/zQPcb4DRjKyDjNW50S1wFLqXhhZCOfaVkveU/AZ1v4AfkX8HZ+XuVGFT1rdNEJr0xxW
fXfDwICxhrSGznRTlNBpLCJR+lD1eLCg/QNgGvOb4DLqvppLdAonIhnmF2CBSYPQr5uuabIQ34gN
GAlXGNHiF2JZdm/AdfXZ6BHIDQ1LvaHiF6JAEYujBpdTtmZjk8zWwdKcHAv/Qn90tJXPU9ucJb2V
/G7HH8zyG1Wt4qeMXXeegxQZDpEtNtPIqzx/b9Jd6NBFbOm89mMhUZ7XQdauWHy9cNTDNlhoS6IF
jfmMQUYAo+YnP0ZQtFKMVbCUWoxg1vv5IaocpWjjibfev0lvEnMGcpQqaAKFsBsJod/hnf+EKZJv
Iut6nE7CodgfOcmX0GFpeKbqkd3TzKxnK9ZRml5StbmhWXQLL5OGbHXn/d2N4UNBAga+6hFLrNR+
s1zF+R5pOWdz/+gubWLaDbvv8Nx3dK4PnfsB3VWESnI9WnWQtkaXFR6aG+b4nvG5isv1pUgHTNkz
J5RlQ0DDz01SL6fPeg26Io3IXhP6BwjTBsijYePgjSPtxsEHiiiigjFgmWBI1+2ElKbWHMRmS7Ww
m+FIvbnVf7DC8Ab8jkfBUZXtJb8wsxxYGnLbHmZz1FAAYy6H67uz0owUas3J76ZTL+IHdsobyvRe
hpsjYp3NG1X9KDFpRt5Bn6XrL/nuudWXRgYDxEUDK2y//pZF3GFbdP4dRk7TWg6FftVpe0xEo/8V
6OyB2+nhttMBU4tisrPPU3rCw0bkakcAhJ8VzspA890mMg5dAXsV2s4f8XUoJ3j5YLd862pp1xjD
PdYuNQ4+hfwcYTN9bAgjwuu0E5x3aat8A7ZK5bmggtbpY615Fwk4XdsmlpxA+oaDiaIlGWGBTBt8
hl8Z+QKVD7zXfv/yUXGGdN//N7XxOg8qY16rrxHY6bX1/6TKBEJVHxQm7rjCjCc0kqN7tAx9bCxu
jtoLNIB9SoQizuQqxecc2Uisnlg61AT1puBIsi1qcpWUshV8cHnQMSUwhEarik+lafcU3pujETB0
Rqy6wdgCQC/NzUd5zXgC+vdEgENwNvqTT/R3DuS1Etu/Jxt4h+eaTKbGf1j7lwTcXK+SLIMZ9oxK
S9wW7Fl57ZdsclMJYoHjzTo287y4L/8vKdtOqed205bDCHSmV+HSAVfmRhLkjoLPCl7y+79cYezB
deJgDU4zk+SEiWJLzprHFvRdZF40710hBVKZR6Um+CVGGsa+sazmTp2YtPqiq/RQ5w1RykODEpmb
C0NC2HuSE4sVDEgEJLHzVjqQ1MjcJGI6u/HuLsaYliU4YuR4skw24L5MwPx8kIb1rXLJQluKgNmQ
o8KquY5eK6P8eEVPGz7tZz+PevKj6Utem9hpf1hdEWaEfHrdhr/q8dH91fevZjNOGUvIatDXuJam
Q/SGUcoeJFXvZ40N2oX5PwErobyTlk5JCwBIqx9iIt/AfUGxYgGLjF6nsLXz0G4FerjzIsN/Rx3S
hhaAsSoLwJceKX6oZzvDh29VbRDSb6XkTExBAuZC+VfpAwfpkKwGoNurTlROn6lbAd3OU6l5bK/+
Gg8MkWwoZZHBZdoo3owocD7l23KfyPfCJI6eJCRdO2GDm21Lty3tyDLuhtepQIayTnX4vcq8BTVj
D4Gs6MmHjKZy6AQhCNDv9NXzjSXgLRMGG9WTxdJ1rsFac+FgizdwtFto8DIgygt9VfD77936Pye8
F3cH0d/KhzkwbwPL1kQH0clcc//5z4FTBr1wgQDFG723/bRSqODD3pEpZvo5Yv8w8/qQzrrVsAJG
D2LzdnYzoDpFvFuJB+8UR4y+jTZovPPBKdsuM/xOx6QIPpKX2SNrTg1gBMRPNYk3bwe7pR1upTJM
hTnqncK3mDLYTNhQKM8eBbeKoDQ8Gvmb4vqT2B3PCCu59pGwPucZjPetv3Xh9OPzXDO07bJuncGE
lRqLwa5tPZ1hUT0msmUBqXQigsC6nY+xOTQuQcMkxsdPuXaGUh9YCyAHofmHSeZUpUzu0UQlO4Ev
62uVIV+lrOcYq+NVrEkx2oA3+5TUhfc49/eUmjPcDfTPJ7Io2gaepw7Om6lHWii03ka1CKy4s+b7
0nfnboGKDlSa4yKudxgNT1sy68A5O23eO9eQ8m3oC5uuALT94YSqTQGnnv2vO6w0LT2LOLbBuHWX
la0yBkWR4XEQ2tC3hoXIOxkUpVYrG5iskHzDfudqD+m/Nr03YuE6ixVamkJEqQyCM+EeD+Ti1vyD
vbrN3423iqofQ/NT15yr9xh3YKBGc11kpCag+kaxObiN2QXccnSMYsVsztXafULuyuX1tIYbj8TR
2jcv9ZMFYzgWFvBHSIbx94gxMIUcgh3ZiPsJ1aQqtFPAnCGC7M9Uk1BBQR5JAy8ujnSHWstY49WW
BmbUYmC62RbMQf6/hJSeRAL+O89NwwNOzXYyHXZhxjBstq3THUEDoKVSVuvJJna64Edo1HFf1pDi
pwpTsbhtVNvivSIjSXkz0dD5URcVzmTgbz2LfW8cGeygdMe/KML4TJpSwgXe/qoHVbewFJs3k50T
YleIvAUa782BlMlejmBjGqEjDDsKqfX0pBjn+ZMsQUD8fdVIsfywTxQ5QXHKGsoLxMrg3+lD6s52
rVNtvTRskJr/faA/mYL/XPfIhh8p7DFr5EM+PJn3iCbdrahLdDBcvQq01D2EODrQVlKB0g8cd+C5
rUMPDo9GS7vrIUdzH0blrhAmXj9kFXCyIXmEW6T1UKX+wctT9qKYrBMeB9hnEWzwgtyAbTzkma/a
kTFLCplT12PpjFZ2bM4LunNEieplU9KjeJqhz7KJZbUFwJQpWvWSHHr7G5EhgyIIN//yWQ3yVPhN
Sodmm7EDOLJvYkqklaL8hLCTxvxgLCDu49d8wCSdywQ1Qj7GuQ+qDVqlZo6G1Ai+vfS0sYbmFH5p
3e72Qv41yq4PBbUbNU1eyiWbIe2m9QEahZ1rpIZSxOocLs1e3zqvczt/5oqpYecjPT1AymKwhEaq
pCikYqTTUAmj/0z3d4uYC+hnF6Mw5WjSPmB4/+a9hPF2dOdLhuiqDiu0hwMhRKFu60p/VyUIEpUZ
KccG3KbEJBWUuFT/5Z2Uo8CEm29XJwk9oRZfISb9gDkV/C9GdsGWVs0q/v9QczKkrKNNV8Q7aKMZ
P1io4oewyFSZbfIdBmfAoSiiTzK3Z7y5XIUr8G4RjQyGO12mnkxPBaUJkf6/ueZbVG5fi5ymYdfK
7X+ubxNTqwd2QZdrQfuf2iB1G/t9lIJ+VRDKBKPQ04JweV0PHQHZkijfmOF4yysdqFjtUFnBqK3Z
CDYS1P3ux4DPzCMPDfB7h5gMLxElcvWxzsu0wlH087tB7G0EwNPHHfU4vp0YNJJdeMEpH8sVXjdQ
OsPE2WZVFGJzJOgIwJ8AneXTaouE6V4ynEsK//Hg9mmG4DPjmicSI35RRelhHPAyyi7z71zYAzI8
Gxoxnzv5ml9eVnog9QI9dgcCr67pq9r7tsh9oJiDEBQYXFA1d7Ojba8vJgbZh53B9sKZGrPZ8Q5C
Rb+s+ODKJT68I7O9fRi+naYavQ8MW1B6LSE73YaeiNL9aHLcGQ1z16iaZPTDZeRZvz23R2gacDMI
5kCWt1hrM0h5aNwVcsl+4t1Kj3zmiB9Sd2vKXx+zT9ClTfG8Xo1e+zItx/FwMDTmgqWQPXpg6dLv
+9OPwen+/FVqJJiLiLItsg+T0ekdV6Ay4BuxNZqq/Q2a/l22GMGu/4jRicgO21dIEjddVWNranCu
96yN/C1Hcif3PQLI/lZyjwnjuVNvIdd4KzeVnJXZOZnlE3rgOUDo4Vt3hVnX5I0W3svITKX/qLUk
5w2+VJsgmT9f72MsLMcXCCsroXprc1qFVpqMKMStEQVVvSv7lwzkPEC7efaHVd65VtYbvi5HMau0
KzYbfuqufZUBrlc29ntLPfRXNPfDmOt6VN9pIHIFbvTOhJtyjwaNQyMPdWCces9VkCs37qhkmGRc
z9TbUKwUnIGhevGGEiFOHnQAq8CJsBXV+6X47xmumrSVodcUCqTuJGTJFVEU4df5H4KA6uUgU1cp
tn7iAB4lQ8RtIFoLKPtY9PcdHg3Ym/9VW4x5mrAXPsUwWCZGfMccHZRBBTS+vT6e8IZElKQBXois
8bEz9VH87ZrVa7G60j6SY/hZ/M+7A5+FBgnzNM0RBygt6KF64rWwGzy5nl6mEcUDOW6JAaCBmcsV
Ob3Td1xsGpFeAzgXmxNt7NzWcwjdSMwX433hXFn/G0VVb/8nr3oKJchCfQ52/bQviJ7RF9Zk+Jx0
nOv/vPyaGlqHhqHW1nPwQP7CeB6sbe3MErIYqNjJKV36Zy96qcvBMk3p+4c7fBTpec9RlaalVorG
eGWHP1epcYWjjhskKwRqQNbnLhabmHhyNR3IXR3lX8PHr1VByFji6U78AIZbxUwpZtxy/NrtzHPx
tM9e+2/NL8nDdzek4mKXktTs0qqzedcCMR7yOlIe2cGcbNltM4HoT2BT/3ZgBsxZeRnbM83jQ9Pb
H96BHmqqfIrcZWjQdWT5nCeV6I63+dw6iXA1S4vS/c3UnLFcKYILov2t3HvPnwAbhEZqZ3IE4xnO
w6ItLvNEL4dS2sYkJdGvvqqothL892axAi7jhjMBd8quHnntwaa7sSF1orRRbS1D4E9kAXTfybqG
kOKBa0DIsnOJfbtBwY7KVdfOIWs5ooWifHVcs/mUsIN55crT/gWdPG5nnAOe1m2zB5+Luczzjt8m
+mkGNjnBxwXPmg+fqYGoj4eTy3sEOf3h3H4Q1pAovllk/YSyylLql98zl7cDOmJJu2KupRxKekbU
gEtr0CA6iFRQyVC9fVo0Hjf9/I+D8RNj1bqtbKLgr8YqbgrP7F3JnMhelr4uET8WM1RSa4FljdyF
c/M6tn8fV0B7/v6uR/hDmg6YIp4BwzQqGf4db3SsokqfA6Qi0/E4u7xxIaHNDDpDPFKzpXZggF6X
FJCWoTza1jCyw/FhqbdS/TH8+6U5j1inugszuHgL4NAcV0b3jRmb0BYGou/P6drusyIWPmWLDd0o
e6EzV6mF2pMJe4I1zhFZzMUvI5M0N9aZ4z7qC58E3bqzd6Mt9s7wxeGnjV6g/TIGe+MfliNoTJPr
6i6IS4NHz9qLQ/+vZ56anHuF03YhvDqyufgvcMMNp6LsNqg5x3mqF/5mYM2tlMAaZsxKOTqWzcSV
lGO+Uzr0UfYsHPnvyx4POFghQOE/U7LYNn4DMhD0f4sld5pYE3PbREWQ/HDOQA4mF5gFtFIwj83r
s3YFgLff0fNetHmpczZrF2JUOkMWtYB9RBmPPthf0npy6bDUoi6CkAR6aPzcl6O3lTfZXFvTRu/8
fWzP6GlMonNg8tOKOCbVDxL/aU6j76VTymtVb92Elm9zfRjgljSCi+6ngbiMWqsovmV+R72c9q3S
dHulgCdDrXgY+BBo8KsTMyY/Xj6zp8dYYIoV+UIA3VkFtQ3stHnRuiKhGNVHobRK7VjcB3dNnU9Z
t9jeaCYomuLEOtITn1wxrWqlKgnd30rFFDXaHRDRxr0KIrst7awDD9AbeCPVZw1CBArcT6VrdnR8
4d4qoykraXaiXFqJKm49zVSc4js3/kFdgb4HEjZdhqrK5sdYI9+HplRJfjNKzGeWtx8GjA/uOp/o
/s3zfUieZKX8F8LtaW3CZZCVRcjkip0Yjbhhx7O5hzF53FD84/mOMpIZWsa0BuoKOc5gEc7JURjJ
wlXv39RdwGckhTRX0Myi1lS6ytcPuuQ4YlU1wKUdaKULEoKy2s3ziW8xldt+dl/7eDw6TKV20Ytg
ysyKNKmXbP3/ZgZW1NBP1e6HrUBDlFMhmcTnEzTS6PtX6bXLNUuzT7GXI4YKTnn9XYejrOluKK+3
K/B6thSpT6cysIQABU/Rou2Ww+c9TRTB8vbL/A9ze5zrsvAcF8eKR57tS+dplrGa0BcgBDObZakq
0W+jfzroJEnBshX/n31T4rKOKWnUaZ2neuKrUH08J38Bf1l2u0cPVvZQhzUXHpZJJf3u0/Ks6Kdg
8FHdgdrs32Vzc8Yutkg23zqskqdpfsep7VuzLs0+6B/Ti19nQJzjo5p2ZU3EUTiN4uFciX6+ihpR
QDtP0coWri5klaivQJqRyp0rt2LFxn5Q0LXLaHrNNlkaCvzkny06ur74ZMINIj2WigNG7L+7DQ0X
Y4TgEJKUY1TV4igXhxNo0ziipw2oU3KiXaMd2COcOBGmhciEN4HKipt+irygFAUrMVmvFNVE6lcY
T+2w9MyO8bpNEXcdVGb7xJ0Ahcus86qVEs2QBETG5sfxS1GoPNAOzo3AwF+9ebbweLBalUX+Q90C
OVccE1M8Y9S2zjsFghz+CA1sARQPFSA7AHPnjDFKlM4x3BswdXCf8Nvf1HrgJtdgkAiiu6N572b5
DlBNWgnzCLp7lGeYPzX4fuxv+96EgbE8Er6PhybZ90uPsKIEh2+dEXIBh8buYNPGVuvWIvc/+4b6
W/mc73eVIwcv+Xk99CwocIjuYTNot3e57z9qb1ztwmLJORMLU2Arzv/jr4P2RDD4Eb/f363thBkA
WsnQRIoWWAcQsrq1e+NKgRNOuQM94Mwi2iC+ifo69ctYB2alLXxRuaOF7xR41r3/DhH/GgyyzLFx
7C9N6S27JOSzvFwvrhTWz9NQmJHJXiETvon1GrVLnBGe/DpbBg2wx79C57g9+cR54I13X7cDAm0k
IAUu8+3m9ctVwXBKYzQs8Yk2hweITxGY+hVsvIWlCAY9Mm0hDcvsXmKby2lEXGLy8zPLLjaeTHOO
G0ZBEUwT3DOlk524qHqYdN7NaOGje7yh7xU1C1NCBeoYsT9soWfcLzObKUhWpdZ/Lt5//8HqZl56
y3BORhssjdSx8Um/jm3oBRtTYae5sk2LgVY8vLvRAaBksVyxH5cNkPTv84r9KhZLdr2d0DxWKsJF
P2PxwJ1coc/GQ8L8eOput8qS2U0hFGGtfShsTQ8jJylyLiDPPLf4ujm3Dl9b99ivwjqVzkBWcPFa
1LGUujMjxK1FiazGvBudUS0OpRt+TPJWv11E3ZERLtSqeiWbC8VljmEpl182+fyqz/Gl3FwLM7QF
ugS6xg67F/zVZ7kXuZ7neiEcA+89PkM4S5ulDaaJsWVVNijwMa344rSFtJmqvxA5J1/Gw9csJcBA
bvUGTuDU+Fc6TuAWb7+Mt/qM6o2AUh4i+uvszjSs9Hoj3da1RJd+AOayvZFAVrUJsEEIikYYIz33
AwSMKJ+8ShJOI9ZF6QzQY7dswBnLI32VbW8B1DD/ActuASxBPLC/HY2+YxK5lDX+olfzJm6CZkJR
nYfvJIZIJOLI8TRB8XcR+nAiE9Iz9UJ8hXDivpyr6BTOSYB2Z5Fh6PH/z3084SB1ghxkDTeVOM5/
4+tNOxYXDhPoatyxJFKSNCV55ejhqnIbsXeEcJLJcAscScbUfzTfUsHt4TiXVngiGHVNKp8Ra/C+
u5U89B+i+8AqzbElWlsHNvOa94EoIEUMilchBQbyCxuUoKrkyOqROUQfqe3bzfDPOnpJUFX/73cR
tc/BtxaijEMWXY2TePlJ7x7nZBYMSRWen3B98OMFQuPAr6j8CaCyIQj0SJx70JOUJXPytxNjXob2
j8aLTnCXfeNxi9aF/9a4JcEDyrqMaRcOzGHT9FVv8uHZQLz+QZ3LFylDsjbVR0EVcjd1hAnI4OUq
DdhORt0Gmd1jCscnJa1TQ3eWsSGZ4bCi5gD1/B5b06DmyV+fjAgYJnELnOaPOLOb6gbUERUTnG3k
J/qrUs/akyXkIW/QbgAuzRXlMZEK/HEGd2DHRWCvJ7sj9js/x3otxy0c8PunhywzKRjcJ3FOMQ7S
l5E6AO9a/ekzzPclrcwAMnfGfF71ebvci3IjisS47x4rQh1bds5bv7jmG50be9MyuNuQVgV6L/cs
NH4czdZKYVv8aAjwwJVQ1jaDz7tRHcOElQeF9kgtFOgZFGtSflaqIkuXTLL/VA7y4QkwoKCOoEjJ
fl85m5FLQo9phJsM7INcZM/Wg23dh2sATPFh55Slz1R9LA8EcACnPy/N8EnujdKGU78mq5+VzvXH
1tQeLY8wznKqpZymE5V/0L6krUGmJTbAOnRhxrgshnWHTVVuLVcosP7Zoyv69VpxwbLELyTTJBAj
cSpoiXVyyl3KGJ3RqxXxZvonIDx16retH5GXRilHdSxV87Er4iQL5SD2rYxZuy6RbIsInipxDcBs
SjuIbCIa2FKQBuAFIGXYTDcD496cC/2oL0emq/EL7olLfj5x0Tu2jvGEG7LwlL0kNFtM+uTNwDuu
f6bz8G0ubgVmua3fh1ysJTP26tl43YXO6JrSs7zNz0Gfvumf5UIFxYwg0lkGpqzesnWXxuCb2ERS
mrsOtfAu+nFMGNLdP93GaXx7OCV031pdzn8L9TUwLDu/dkPPxZ1qdiSqvoce9f1WIK3/dyX64phy
dEIzgc/xDJaJwE8VmhWZloxZIK3gIyG1Zisoh2nU1LciZpQXEZboT/15+x1GOsN9qtE8zSrLDwsG
u/s4Gu7zto4DNanKyGBEI8Vmfuc4pO2lB/P1yuwLHhLuobof//2nUwf8RLXGOLNOePC0ZZYjEo0Y
9M+yv8dlhhfQnNdVoK0l7/0IJOVqwPkoaJLNQfYKu3jlykhdvr+v13g6K1na5PT5OijznFEwn5CT
IIJYSq3K6ShORCME8N/ybu8bfN72bwtqz555lKb1sAYVFsQe3qTYDXmf2LG8+1QzAVtRBZHmvE5v
v8cXWsc7VNBbB+a5kbmc12DiliQCr3YRmsaHH64zCtgWFvdGtrENh2bxuWKC8ELgFXJgX7fOOD7Z
Wr5CYbkO82ZBudbbIi+zZVpgJxtSsoB1ASK8E+rXEvOXzhOLHdzM0VeeWUvHWF47PNlw8J3T2vLh
izH7dXaCCxSyleJJ3Gh/fXrWlFF87WAisL9VQCaEQCwNIUvOVM71qllNik+Tov1ZCLiQuROL4J8G
Muw6owPzVLWLsdcG1BQY2QNwXwfDNfmdOblKbRTmLBXtT3F2MScFtmKAFDh6F4Jki0BFjQdCEJqt
ZpsykXIdAi4ETtRaMC9Cc5idrVWyOGlWpUjrpSRZ/L8dyevvjMhtIDhsXrbJDtjWxunQm1In6XM/
4Jv3s263XkTXzkTuymLHjupMMz1rVul3fXLsx5IdtoWhcZcx4ds78Z0l1WZpmanrVLCd1qDca9f2
RiTL/Ikkoow8b07WvkpzkHwzM7BiiZWa1h7VChATaM8x0d/mbtZ+rcnbl/+XCDeUdnWosc9KjtQi
h02yNXoyo6B/Y64TUCA5J+m+bFF+q5L7PPQtWe6qkqN08WFhrbUIzI+BSs79xFXqx41cFdBh8uUr
g5+4GH53gZayiWDxmezFJXEfRVYVOGK8aSnJrUxzCrEFxsjMilP4PamNyq4Hy+TNMdhGGwO79nCA
qa/ZddMszcEgBBzTl0tl2guRBzs/BzeROVOnCo6EgKkUznMdCGfRmX+QF5TSm+ETRh99XGZIfv2K
CqrvHxlBDIKhlFyHtqwzbCzqGFWzmZirBFOnmy8TyWq5z9s+sQ4ny8AKZXpsRwReuSbSX+f7C/B2
qllMmwL+pypphSlJYmOf8MFoQ52gHApfEu14rHU4Ln0S9Exdp9HTOEt0eyAJwDAwh1SGNgTvOq+h
j4K40SZ60lgsseTlxuSl4Y0uXJH/EFVJ1u2BC/JHOi0etypqJ305nkViOAcLk80txu7M80e/ouWt
fy6ITG/ppitLaiFrVQii7/f3fRQJSSQnmxM2r9g3gqgh/KrWQ96eHQKF2m9QMdFaW1NtBj9OTuiP
nCHQDKZOCz7E4rPtYhSYCLNMpBh8gtEpbZEGbMT0PcsXRo7WFn0kazG12bg0hhUG2FmcxN19l2lu
eJwDF80g56zAGZpehYnThOzUVoZKjeQKwB6k15kzBx38Lr/H03TFbQNEegEPjIDWq3zpPPQGDi0+
v6/xiqqgBFZ4d9UKG0UO0ZO9qT4uMQflb35DoJCRT1EAUi1CbKxdL4KoLDsHRlfw45cQOoqnpLXy
yZCTt7gef2Cg5wY2qW8xaYY89Zk76ap2Kiavry0ebOf5JKqMBT6+lpKf42MliNnUN+/kcyB7C9WI
FkqJh48wc3obl+1PgbbYyjtHUGqWXmHQfntARGwhHL5IiZBsGGrmjSxfD4M1VZtQCeOhA2NtmTtF
o2O3jQY0CXL61VnuoNb+mjhZYboigHtNwtdhuom+xrmPbIOVdDOC+dAHJaUIc7F6vJ4S1FFcfwQd
JrUNQ3qsf8kx5gRhGyuEMQu9huG2g+ZJ3zbGPMXeCdjOiY+z59feyJJEqAA4WOG6Som70sMZcBID
5F1hMYcYnXlBoWpiYF1xUPZFN4uyokZfpwo1SwtcYuBqfSCkC/+hjkJzypxloodkjt7YYke1ziYj
OSjE4s0SQwBF+vn3g/fdZsYxyOrzTuEav0zFODQjM90cScrUolp3rPLFHASmPWPcjLzMpCetqMUa
JdJJ+A+DwxEFT0akk0g1ji0jVpZ4pyahbQD7m1d4r+xwY5pi2YJ89YKjZnAcwpKzYaFyEz6AX5Wr
j7NACDlvhNSg8ilzS/AcwVx9S3EYBZY5WYHzGvUfRonQmewOFm5jaXQ9Ax59vslHLfZq/VpkRYnx
W9IEOCGlwZAGyxaTlYhYPmj7gxq+2e0W+d51PyXpB9OGp/4p2M2tZ2Iemsxc9KfyY6UP8BOg+04x
7Aig/n9sEGnajKtrw7BxMvfhCySmmQd3s6xGtaw/ss1TjgORymU+ks6dg0gALAaz/UBWX1VRzCHc
9dVL5nRZmyeh7S6bMQ74t1N5bTBTqFbQMkpj62Hbd9hZKy9k2a3vYDBqJWqN+U6yIzWo1V+SFS9A
NHrHtoVERxrvg4raw+xx3UvC911Q0GyJzpnqgsPFUgVUPM5lYfw32vxPLUVNR3rIidbjVBLsFkBT
EXbb4nCTJuCZzB1XwJikpA2lnyMBgjZu7CncOTyJWA0p798SYD9/kuZ4BQShp4Ho4PkCB+UuXpWK
Rv/LZBDIlSOXz0vSWyDnS3/ZzW+Dy7dIelil0J4gFV+huE/BXw29b5W2Vqp+LZG/c1ntLICe+BDD
lqSvYqTFDtdFFZeGqzTKvwTLJGX13ZLveKPPNy03tQTweajlxyMp2zUnkcdHFnDGJCmLI9GmoT5L
sFDU1bHnq6I4M19ZRrwL6ckF6rsdg6htPV13hf5XZWTIdHVhP5WAga01P1IJx0Wu5lrLVZ98e6oW
2EUQhmxe9h68TOjiMcNEMf/b5UuPTS9DvId1zB5rWZcIOkPdcHN5BoqkMKFTB0/UVjFMzhC7nlbC
YS7YvhGGOKTec8yBf8KXLYKyRd13c7frTzZ/VJNeXflwNzmmRJ8Yz31/DAYWOtFpiDyAf5iykSUX
J73Ex5yTkeks6DXgJTAo8y42eI6voJXDks55mlDeEB8fPqH1THsWaCxy6Sb0IvSoXfMFSFLenMRg
JbL5GakSs7xn+fWSgk3es28g7lsEI5IDmwnDaHJnIO68T1Km/F/8rIKHOtG+TgTH6BEJ1n6ypJim
rCNFj/Sr/Jpieb2p82I8vYLBSJP9f8yP6GlEswMu8d95GsQnG1Thq9M3ymo7L13QI+Ynhw3coK3p
1s2zo6PgTmCYss/rbJ9yxBIKPXEtPPSi2iM/u1atvoQJpG3g9w9bvWC4E2VSFVH4OQy0LofSN1Cz
Rg1bWmdSmwO3NDMM63orCI6SEPbF58XWPZxy94P0Bokrf2c8aJZYdW1A5sme0KRL0jeazxkHaxhm
sUUqns+NcaXYFcqgtrIfPOjNEdHC5YClI8KZKsU+1Fn2qCEiKe6VMlyrZNMnqNjgWprtZOeKSxZs
ITPVG1veKNnyuLDVC/KcDgrlKYBOn0VhGxQU0tkfWYgvctRNLqu9ix3zysW3nQ7/JyVfAdusC5Tu
mHYi+jI37JqYbXawckwOC+fg8opGDpHzWhDs5/B6AWN3MLQ0INtCQCGsKDrcR2hMI/0rAdJ4d3RQ
+U5/cIF88ROjejPEcGxQ+m8+fZ/lv2a5CprW+1cgDhc3/XqTv3ViciS6I18MhWaR994Nd8aBeyHE
XZ7lKqIhnc0nd/YbfQs7c4MV1E4hbAtrT/f1QVP18exrVhAQ1cr2yTc5GA0QKhXoufSWMNunTX91
5ZRKR2/osTyhHiP4mrtYnu0/cltD4EpgBO2rp73xS2p4MMxjvR9bVYgweH26u1Wu5sw4yk/uUm0Y
bHfGyBm71IAMi5agYLxXWDMc6KxT4LfbrqoDL8G41nwXGxGJXyBWHY9VK7xdyci2E/HCuJi5Sih2
d287gFEXpmAoEzZ8K4xRVh3LZz2oAfUEoZVSiFxTn2OmsGrHUObBj8ODsQfp//iPldP5O5vocZQA
kuYxLZshpPcxFlQArWpt87FQN7JEn7NWcnny4aMac4c7zdtDzeMx90EIRR6g2ka0Y9fMUqac+mi7
dzmyb28INrz4YuEkkg3Ehvfd0TtFoupGUr8CVUqhfTlx+PkDHMWUTQ+ViBzQ/AaHYuoTvojf0c0V
lEujG6QiRvBzsf2lBBeLrqteKyKaQ2Cm/RnLykIARnEKY447pZMN6RLpFaf1smc56Z9JdAYBaw3a
RP6miRSvd4bPxMgIVHbQlI4+H8ihoSIwZyKuFEk2IsKeYyzj5xywDi3ksDADRxE+AzAXGdRE7PmV
qmmsMSmZaB3gzaz/gCOfYV3EGIPyt+H3qfEx54a9x8eWaqotM9h8xJ5d/gaMu8TclNgR8X/vw3QY
wWQzXFz1vMFwYm0NuLlOfjXcgEMK60z1APUSinrkvrhvU1+4w/SjiC4j11BB73nc+i2yox0d1Sea
9pVyArkJH3/91Zv0d7SuqoKw/TU+chNtbhRhwWz75Pt8qDCUjBbH6O3CAaz7ibgZdhmXxrLqfToE
Pcdi0yMR6h5YPlJSgEHJR+pC/4dZWbclVaL4rpLZ87JqMQWBXOiqujHDxoOXr7LMldxBCWLY1B/Z
uXirdRzDrtN12Lue98WeK8DI9Xf6DDxrWOKmZ0qg/UU9/zjBFW3HHotaSsayNskO+5osmHWYaxvT
7DSEOsJ/Vxk/3AXt5jIK9Briowpyf1w3hGnBKdjVyCKd9hIJA/zlidZePWTsFoYv5wqc3NkoJC49
OMTmAsmXhFThyQmIBx60uPxBZA0gj7yIU5JrTKOui8ev3PGju7gznMh5a5ovj6yqwUx6saC0RFSz
RLy/pvcftv3L8lTA4n/8lR3JViOtT0ulMgSzbVtfqd/689/syMSHgXBwm8A5Jz8AQEe12aQEde0p
Vn32iJQb4mB80AE8/j4OMXU4STMWqSs4eu/Zlh3m26gKSxp6qbHviJXPc+x0xnPFjxsYtl7MFSw5
svzfNstJ1tXGRQYtH2naav1DA6FdyQqv0+8rNPIWmkYhWEuQs4cF/EhihokSYgbNGutQgwpVH5AQ
BIE61664xykqJ2WYukHh0YnJsOd0WUJD+mpDSbW0wTjeKddQC2cnXG845cmkS0B3/HUfwXC4o143
XgFeA+qSVkDLDJBzhbjZhDoTJZtDYHEXTiwCLqgv26AW+GCM8E1bG3+AhUbBzT7k55/POJRbKZVf
CofinFuOyrgMWd9RZndLCoVAyyIODVnNK1gX9VuQC2is41BQlXXuphLV7VNlBi3UlmTSs/v40ccV
aN38m+Ri63OhsvIRzaQU6/pcUsoEqs26G+KJthlObptFNxan7GclcZ1gDMtuEEr4tXBoZXwoUN8N
Y69hkIHxO+t98Dynke6NcOCaV8kctdfYVJJfxpqPaX4pYOIixsaiEASotQsDE2KyN9bQogSgx5Vq
HktAO9XTTPdmzlyPRd6+T24zVX1v0fFuEEO6QCuQRMyOB2bEvD12+U0EGhWQrfcF2dD7yNqbsVCW
k/qj9uqztLArrelGpMXcgeaEbeqesNtU8Z3krs7ALw6h/201uS7QdHFD6LxQsCfvoxfgvz1zcLy4
Tznqy4t4P3MEpb9zV9pg+Kv4VSNLSiQXFMUNiVmLhIijTx52fXBy+xTtP7xkQf24akeVc0dXzE2Y
LIdDQtwHQLLFxc9YZIKFySJtflBX1CbwiHo0KZq5M332TSwODeR0dVDMHh4vJNZSIg/vzfjP+RHw
C7L++KvNOSD2OZcFXQV+3MV3S3r4Yvcs1u3LD0rwPqG8KJj/EtYt9zkCO3sN9SOo0SsutAAcsUcF
sKJzW++Y49hI6JgBZ5vTlG3Dn685Lq4a5jqHcSmNcF7pAiFcBRp35E32zSSnlDgfRIRt+IBvPq1a
Ta8112lsnrglCChOUZb9T7kBXnAnGF3j20+vbAlF4rsKsPA2M/Ee1DRKQtMc7wl7wb/WAZwMxwdF
M96YXh/ZuYZ76VBLPJ9xrljlCj7vtRVHy/L73U+jJwnj2Y4osuwZ19hxhGm8hi6gLJArz+xCWBUa
U4CZ5Yur/P7TwCtLRWtQ0gvduc9LHvSEnZMCVIysKpm/3RASZmA8bEh1kdZ49ksAodSEh9nHggCm
3Vxpmhg0advQxNzJVm7gHSTdzjyKZf7tto/N0JruInONVtAN0prk1n7iT71CPFhWfnotiUh5pY2X
W9xSkQ2UzQm97RHseF0UU1mDI7hTm6aHnUI4ldOfORAvyf/dwehq6LP1U8bsyEs2zfBYHeVvHtZj
QGdrNsUEHF4DodL7hRhoelPym3kat61lOgOTch43l4QOHdSQqL+CV7EyASUYorOs4e/WyquLFb8d
gG6u4h+gxhruLM1T0DQAp0I97gBn2WqG1iurDT3rdA5x6HMq7HMS49Uf49J8IcP0qPk44c63kW/a
CD0Ok0IBbV7HSqQVUBZ4nSdoAfXmgU/2yQxj7FqhC99KVERN4fbOmWGW/qeYxe8Tu9fMRBnWldcd
apQVatCKytfkXgoJ+2uKmCmzRNiCjixbMy+Jdi/ViVPBqXAbVJwPAtcbAWn8M16ePCIOj0EJro4f
JCmaYQIrGyftQ6+xM096CGULurPsINUnTw3jO3QoA42x0dS2MGU0hIzm5BY33ch0n9ZxSGlkHoDI
L+wwrtrR9pRiXZInwG94e6A6rHHnKktAYZIngWMyVeS1+mOhmBFjDRETHlvOeHbeGc/mICeaZ7Op
f0eipHYkI2GaRr48mPB35OM6AUQNz6iSv+1vh/H29GXib9a8F63ijorrTLhnFgn8qrjpZRne1BXP
matK05Ls3cZYx/LXpimLZ0t83cAgmOGSAGUktRRSaA+tHlBVwIghiZeLBZGt334GWrsL51dyvaRg
wBjDVDQGoe8MpH9YudSOHzp3JRR2f9KwO7wNjAhDj+m+POK+9G8AkF7T93/k8FWiJBwRg9UN1z+a
JMxX7yoThXHBmeI3mPKHJF87R2rN2duzER/NQqqF+dbhZ2J9Pod0QjU2U2QibeJAyzdDNQlQdC1t
UuWeeJFrLrlzC5BOLK63XEjV+Bwmf5WN7styM4/ocIhP4X4CHaoxa3Hi+VKB+4uYj6oIVs9agVsL
1rkxi6z+M03P+szqjhfAuQ3c6/su7pg7tRcQpGCwD7PiY3w2HUN11KjQRNra+X2kIEV/lv+0086/
1JMvceJ0ZYPnnHaw7FtMXtt/4gA4XDixR/597KA/mU51RVSUIMyz7GU9lr1e81mfWhMUnn6N2pur
TM4iVM2c1gFyKaJU8EUmiqm0HfWdN6/0Isun1UuOmxZfwEZ5xx5sWPgSmFuvaxWq3qXNhh931eP8
cOZluxvED98ObotL/4z3gbnoVV6d/hh1YeNZH8JQCsLMtES95ol208RQXCLZG1beekl8ZafPQKI2
3iZy/zjJ429kgQezHQRd4FdTbOuiiibCBSlSzxSTh/rYhr/9VZluJ/9ls9Y596keQNpNSU0Q68nr
UA++o4s87K/GQjf5j8HCU1n+XD1NetUrD8L7f7g2xxwP5tkOCOf3zf0Bn4ouZzbCSnSJE5PQW/Mt
iAWQq/01iiqkIWuWiuAG798ERIQQQiaskUqL0opgUYlTyLrcpsBkTwtgODvdgfMNL8z43vfqV9aS
7Kox+4H1asQGzV9nm4wbtpHHzzY67mtGTjuwiEU+ZgP6d1O71a8B04S2CzUAr4I4SfhCHv28AvJg
eZBkM9hLRJMMef88CZEh8fEWUkQ5hDt3DAZpzhiBHO7wTkc+7c2rUJ4+KqtZGJyGPJFAMcxxQqGY
fMXvvgS2CmwMYtgySibMb5aBcZIkgRZ1Q405XQGoZeyYQIzrE+vrA1suYRY5jYLYroG3qJc6HUge
o4rCybPnNTyd8yodk79fYwB9ZDg7wihxugnPgylfMxKoMpv8j5mm4LUxuHY5ZqU5jbQFG3Z7Qow7
Y2QzyBxTG+/kkU5vJa7hSVQdwHDOzU19h9pjNJtewGsgx/BrNMToUlRzsZ7EVnNhUlya2F3XHu9z
wvi7ko35aLY5TTPPuwRb3bKc2xuhN0ipqEbh922rhIe1Vl5APz7wYr8UbBbN5sJjbM9UsnDq4Oae
zL2V810e1sGydJO+JRK7p42kCCkysWdX6d5zCWjeMRQKXyArOre/YGjJDkoMe9R87bYGlh8P0ehb
6ryPV9vBPlo/IiGS6aPjKN5kz9a7RJQUE7ucIPvYtEax4Qv2mv1Z68zQy8WzCsaIFnN3Ud7fWl+e
q7NA1bAKrgnfwkt2T6uwps/z3cy9koUndBMg58rmyNX5mTJfF3VLc86zHYYbrl/GzxFysHGPNQRA
JGShpW1viPkGmXGUMVV+zOC0YShA47r5kGdFWovzCFJh3+JSjLMm4RohvmvqQ2kQiytyQyBps+AZ
W2oS50iUzD9i0OCI4o6p3zSU/FnOb3XCli/yOYtkM/d+U4+9QodWmVD/Oe/KjJPu7kGtvYLLRjCY
kW4xoGhMRD//jiSy/AlzJpAqyT/tr+XoJCNZg4NYkavAWovpwrDFyMUXK1KMDApHbOyBJo3zpqM8
WoI5nRYpYMD9ACSqKkOoMkVI+EiC7yTaWbo/ZpnMU8C2L1SbTkwVs73eOI2Hf9E9plv2AYAo84N9
kEyr4p2ibJWebE9y6OUL+JnqVbpAbFYiCwSUWs1G4TY3OGOBV1zYDeon1athmYTkkjLSCAKnxh+U
5LtMYX7MU4fiGIqh+zXPAdHX+iLITSRWmttemBzbF6BYAfhDduoq0hCBkcpYJKblHrfV46+pimvG
Hk8G6A9y0kNZI4zBr4KlLrXHCs8REfYxFuEU6rpPtvyIV9q84X4XxzuPioiumbaPtlIqo82kz2Pd
8qkVDFXJMzzFXWaGv0Q6WfuHFCHxG4L1Ra8+QvvI0CNzzG7DOB9mTF73nNj+h4aghgUQEgzIl0YL
C4f5E2Sv+xvjJQQ8yAm2tQoGjeFQ7fNUDuzg3Ezu5qPXNLnXlmmk2rUT6Xe7noPyxYnQhr+1qteu
HfGNxr6YjOPC3VQ/Q0iSMvhq2quZz8zPSBXuItgAASA8j6qhLFpl0rZjvlga82ypeMX93QcF5xiL
XajRoFFCJMsS/TJUjTegPetrs0J1yOnoNnBH6lbFqrxS2ZPuAxy0qCXuZV9TN9CwA7zWPpXFjg5o
FxP56wIhRmw+HKMg4AdF4yYKcB4EfgR82n+JOhyk/nEsLtpjnPkVls6NeXmO8F2seU5lvHIS08gQ
8PG4tOs+ym3UfGwhGYPIDZjZNOfkDi2AMYemKe9GlwdQY/7PJH6C7ZVlqsq+NP5ASjMAx8pkR6NB
3SwPg7P+DBBDDfFhiNRldBvYB37gbXYb01q8UVhUeXtbt3szr8t1A2EqkZM2ObcWFb1fXa0wXnA2
Dw7EL0EhuwU6K4ft0NRVEtDT7CC9OFffJb+PhTljNidx4q6Z+X3uVQxiEitTf4CiuYvmrQKvEFQB
bDnDYiUYT2nwi434habktgVfhtdOWECphqk+VWnrg2hWhvMGHnTBdcfe3IFO4XZhMGzpbjKtJcvW
u0iBnWAVoOgEFbCwXIe98PhMmIhGC1v8K6c8L9DrWowBQPrd0iFXsm4u1N+2cqy0ViCPPK3b6M8f
jbMEIAc87GTOPj7z3cbcok1Tw5e3TMiyk30oZFaFTwRYhzx8lqwuO4Rx4MoVm1TDsg3CNE8UjTGR
q5rwHmLEZpxr1YGAqpZRy5dfLCqKuFyAztZhiuW9GJHaNsGUMYnFRnyDSIqg83lpLhic1Wmuc1xK
Usb38DNtdtZ4937m2MIGyaAGyavtOryZCwk1+5Q+PHtZfMjXiQdHlbe8b6xJoMLmgIzGtVO6898I
nOyQXGnjEXilLhFFXOi1w4CKoqdRoCATmGcDDdOY6xG+QuVM2Y1W+G8mU8JZdiqoVnnpBqnWtSCc
xuyQEDHI/Ouww93hWIK8jvcCTsxImA+rVqMgthCEoJM4X3k5N73jNhcELiVdbg9rjGATjaid1tFY
UZAiKxgdfjhPWagtoBCtlmGWjAbc8MyOc0cd12qqeBlJcanIJEh22oho2t2lz4v/QEjPHB99bD0g
A39GVfgYfnV37OzT+o4HDCwopou7wWJNt/5q6cr4CqKWbcLhHkEFX+MSOAajpd2J4IXwsKYx4JCy
I6pgPTCsu0ZfBlyTd7QeEVDI7MLh/SHi0xhjbuFyOCOSYH/kaSTwueQmkI9dtPOfORqYZiBZCBhg
RfYS87+yy+3WedoH6rxRm/fI/OoOmajSts/2cCWojYuJk0ADJDV5hLEmZDTqXmjcZeQ9FIG143w9
mAoYDZGIccyc6YVr1oMSSLxRyrqgM6MExZm4/76CNLOgdKEfGv6K7ssQcMhnNDJguIkIYoqFxBcl
tGyK1wQ4hcK13nsQRgm8LzYvFA+HIL0xG2EN/2o9WVZTEJvwTOpo7ftBhl5HXIiZ6iFEkfp5iBqj
AeNFBrxJNbxPPSrvnCsJNeXVWDlQRAbxRuSibjiRdw/KDXTX1muQLUmEXpbDSKB0e3XbSLKVLE90
t2QWmRSVbVj0UGM66YUqjVwS7b4+gGc5behvrS8RDZpb6Mk615BntQWK3L3+N7zlHGbvBsGpeebE
zQwKPFTx8ALpzgOV+HS/hz2p5iqB0PmqJy9Lva18WaHZR12ElTOXh5qpPprFGBIWDbcWg/+d2AJd
4SYmUnIE6NhNjPiaxN9oBUJprWz+PGhNpcFsG0NQG2b9T/dPSiANU7sY+hdGsoSWrqe3NObdf7Tz
NrYVht2331bcPo/hAiuGNQYbtlBQR1SFZkcbpOijm36T+9ixzfQLhRIpJEbqPZcodiSfJ47+QJiJ
POV0u92bS4X3tfHFMiArS38Md3iAmHLF9mXv4LO3iQmtH8/W4bzlqnqspFGQXKOSKeuD+gavMEZU
/wuvvh1PYBb4v3zb2Rh7BJFimgHZMRnB16+aJuBCLqDqJNqvcdqn/7z4uQfVlmwwnU8k5hCHnoku
ZaX3koYp6oUQ2fuHBTniCvjOMfPx01Sze6JIk/mElhFOs+W5vMZTL+K+ShuQbn40WJFsWVIHq/gO
dw/f/81OGRVyrbQFJfmhJwAl9j5AljdvcDKjxezv7fOi/m5sYK8tg/mD0HNXFAkoIyzo792b69TT
LvQqFh+5td7QLL4jKfAHt25CCm6i3ZzOFDqOXamii0GjwdXpu5DcdDYUhaxlkA/cUlCtdM6l1c5f
+1/Ar/hRxXnnzTBJEix6JeeRrkqQzAtle9dMXxYW2pMAg7tLfRV9atSJGTW6u+2wR5LcwLu+m+yh
BzgoISljwaJYj8q9Yq8hm9oCIXi+wB0kvl/41XN+IqUlNW0+dCW0PEBppqR8b2VCjNSsSbn4b6Hg
RcANc+M3pQQLhhLTUYPMnaIkWqvCavPzZLCDn5vKCOt/E+cnArOyPyqfKA4CwMtmL04yuxXfraEA
RYFGFmAbFFt4I1gMWrbFvPwKYUaHFo2UNjp9D6WFrIZ69/UKHx4anixMOyJGUjef1M0f8GiUHFS3
fVFdnWHC7eWzTcclaDSnVfr/+N+oUHm9pqzA/ov/QlVVXo9lceSYD+zLCqCoTd4bclbxgd9hRLgb
jToXP8F4nzLcnWgGP5raw5BtvocMLz5KuoYEHFnoNkiMDic3dMKoZP5wXIke/05mjKpkB/C2jair
k3/kB9Zm8v4glB5qSkykhiYD1KSUMrz1X39FybYLgCsBjD6h/06TvBW9mtDLPINUQfVpLvAEoA/n
XDCfgOWg/Jd6A9J1Ng0gt3uki8Ohq4XWyidtqzRTkeCQ91Aa8zJGcJX0Cuqt+o4UzmsXH0OT8YBr
0y0NILRRr1HG27PbTAb2gTw6Dwnolfpu33YLZEvBbJCuo3+Cwg5CW72pJ1ceGiFDnAJ/1sgWDCyH
Ri18VTlAHmF0rl+6rE1jhOPXY8YgSoIF8FsOUa5z5/Gj2+tQfaOpDGtquaYkUsv8VDdWHKUiev4+
Kb7f1H4vC5k2F/wDJnXb9Oxr6oYb8C04LxSSCfoJ3I57UjW0bSlwTO216SuF2NfdeGeW0YaY82eZ
hvOrJG+swDmOZVxt6Nwqq4YD7WJaMJo3tVBolbhlUHbgZH/f268N9WKTMf6CyY/xxcjS0yI5UHVq
55+okO8qo1HvuCFEzwFdhquI+Mr9M0zul1ZlZRRLLQvqyBh/grKK4R8VEClGWkHp5jKvBs/10iQW
WWPLVOPn9AZJfzdBKzEM4/XNyYw1VoZj1HqjNzk0SUt+muBE+3a06x07G4qgvLGOmdclzGtIo5Ay
LaD6bujBW1IpwNyv/26HUe16KtWt0qMYFuvmvdBnVyVEouxwX7PdFiOM5zMbBeGh7eEeaFhbrAfm
XeGS48nePOvqImUXOdW01LXVBtAMkTsruKx523hHvdqscchRXuwXVzkMCPi6ctrMNa0rYE1bB4Ak
ZUJvsn+4VHO1k5ybFgpvz2evXG5p/bRxU5rJFIvLNOrmFtlRhFdq7oWzdaqNM96SJ46op0J8rlsV
zq4srpiw4R/8L08D21JxFe8rBM/jTdw5/K6K5wcLlmYtfynuaVAvFkH/4pOJVcJpNJTBCSYIlL+m
5yDS7dJYHKluopIsUJwAnS0rqA8n1zy88lfW+ANDtZjPh7eTK8Fc2AMGQUJTxoRYhJt7MGnWqNZN
YLgdBVkM9zMjAIdMQywItt8s8Zv8ScRyKRkz2OL3sehRQhNtgjfNuPVDPJR2Dewvx05T6iCFwyBb
1LOEc2nToYQw26a5oK8Pycz6FHynE30QuU1CiaQrMcnaTI1XrmTBcqZWJboAiBpWL1SDO0qZ3wjx
fsJxMQmBUAl7BX0lrjgEpYxNhhFOqjpUKd0YxoSXJSNKRndN29zrsYqfVdhntjrctaQefYan5TCT
zjaM96gYIPtm7G3yXT1WLEYKm4K0ZAptPdail2RYMSMmkBLmh1WgRrZdVqMm3+uym3UUQrjLQdHv
SblRINN0chWua3kugUxzL838OTaaW0lTkBN+eHq1U0M3O6jUKij74i66F0bH3+RVQadq3bTXKmgu
sa+kl6LVGDfBRZCqSXs7LP9YG6g4FcBm7PnLPLdDrl26FzCx4yfZrz/B6deyDMtvtOUVOB9DOuaj
7FGqxlM4tWhmIBOjR1pRjONYhTvqBwJkBPKcrexx+k8aO5GUxsjig+TR6fm0SNAx9urhTuPaDA9I
Pr+V0ehFJ3atSyS7IOUvG+F0+fk79zPBZfrZGkNiDBM2VO/e4JLgdDqTkFcEX8QyEtuUZpAtS+Nk
eXxgJ2KMWzcJReuDUtfbF1oPts6opN1VDe9wRari89lgXmrDY787kspLQdD8XFIVGJEafE95J2Rh
/qUNjrFkThNyGB/aCDj9wZiPHTxWPqyq36k+vK/Hu0EDJ40pV+J/Q1oJB3NbZnbsb89hfmiO15oO
Jsz8RE6OML0z9415+178CcCDZaTXi4sfhQvAqjZIyOChfBGBiZ7nKEace4LZ/6j3TzrLB8ABeugi
ZfajDHI/KQ7LTfNFwS0CWjoDGVPSkicJeF5EitW93olvAZfpL7SXX1w90+cXLqCXKaPshotHbYJI
ObX2hHSEGPweMbtswI8jU9ve4Ufu0oLU1/hRL4haEIdwt1s/A2GIn15lleYe7MQi96Ps8ecmXG2s
Kq/DorcjFUMEb16sVhK5xm5ZNxHxe04WTn1QOqvnqKkWGLTTtB3/LV1A0UoA4QgSGc36h5qcJmMD
UZwvM2XpwCa30GCEfupel+VG/PoBBwu5kNoqRb2guwENko0fhCdwqAWNjjDIji+HL5H8ahSc6N5s
P1ba4k1Sd5rwtjM+g3F5Mrpg+mbnSYGgMJ2xeA9UDHI5ZDgFISKFIriQZ1ylsGJGINpfCJrSfmX0
K6uGHPOsmsT2uQ4+yOwrP/PlqxKZf8vG89Di7ZYaF/WWASQl40vf3F/WZCt+agwh6TsCy6A3M/qY
GzCUSi6Y1IpvfMqo35mfJ2PYVL7kB/As8dsnommGsB8Qt/GWEqayFAyOPHuBpVlbL+skYH4+mutz
7Jnwc9+FbOgKgkz/MqqB3Te1yYugWO5aZ8EPr6cnWSvgAmn3p8yH7Mthq/fCgXeoJO6aibXyiTPW
cXRoAdYeQITQ5zdqUDM6nJLXql4VHQ7XhLC4R8mKzsDjq8xFEOg3GFoJa5boCw6IGXwYFch+Bu7W
dHoIbh+D8BvI7NyoWNQL0GlRoUeA0ESgZOSSC7KlQ6KCODskkcP+Sjw2tvwOKopLT3N0pbqm8BiP
CW60P0S5IiuyJeIsQIC4OIm7Di49lPNVVBWkSFJmxDuR1gmt4NB6NjQIHDdg9BPXgq0aDj8CYvo2
anHtRXZuTejaaLaJBVwxLE4/pGAFCdzZb5jmDOG3HB2JnJ5KyxbxbG6PAFeSxMKWJs32bsk6uGD7
dribRe6UDw/5sYyJ7M/ypzOLIApAdRdme3SV/q6ChMNPM+a4Q4e+Zmqhqkx3A8e8BFymY+87+YTu
i0LOT1Qo7qIEMeb5OSZAXiRa551vQ29Q+g2JP8+bxf/Ij0K+Wha5y7rGSwHrJnyGGzFvFyXDfPiE
k0kQSlPVBTKyvAlvAyfP7/8b3/2dOFZ/TQZ7towCFu3Sym+UGZoDnyVAlbidfCJWh1L8p98B1XWT
+n3E/MaHFKTA78U/KngjykDngr3w1Yt3AOe85nBpxtpebtm7mILEPJ3kMteIrwSQADrei/kw9Ep2
MPTkYeQV2yQ0vdUkM/SzLQcuoDKgV0tQdRHEOwzbD2nCfuWx+cAI8Pli9E14FR1wKTI3msYs/mgx
xYygmZr8JxurnzyKDS02SvWs+PKaT9VyFD+qeSXUboMmSOte6b87oiN/YJ2TnVS9WkNtmYvbEITG
gU2pTnDk//gjEMclh0k/DW32gnyzHfDxk7kKd2ltLbOON1xfjNdxbKDRm6wJIkZ1yfTcDSOFXfsG
KmCcKKyYhJJ42od+zx2aKWn+0hx4jAC1WsTb8Dc9kZznuFm4lkvwQmn4gYWucVk3IQc96caPeUKt
Xb/3T8ODMCfXxUBL2vb1XoVOte9OWTnFGizNbchj2XoPx/rndbFDVitbimKqTAtBF7xKtnPOTAMv
q+I2enRn1hOn8qGxU6SJ2XFvMAI3lM+EYSMznL0Q+mUJH9995KB5XdluXOyky/q/dm4bl/PcmYkJ
ViwVzV9o44mf1ly0ImrEbNFHbvwWsP9CF343eEanmezzee/US4cJBpc2Yh1roa04bVdZb6EbHdIH
LUj990RgNWs0XXIX2WV606NVlaG9vsWC9mBHQPpPJoIfNUY+OqP4cHl7Ha7KVIn+QW9U4VHckgg+
HaezA6Y6X+VeUKLjpNDWGa13wJgxcn/kt+FOXHe6H+494+L4K5uizvM7J0RQoYvIr0Gh15TCG9yW
5G0NMpSmWoyURR/64isZznqgqBmfumIVoXgPkkqpr/gebVIb8o7nVdWStHM8fc5rY5HbWjgLP6Ob
rETLVg8xKe8Aws/Q4Cf/BIk6jbehsHvpI/qQ/2q8/AvZq6VxqHXICEAObYdf6dqYKe2UtmNG/N7T
wbGOidRy76AwTz8y0ENLBQDvd+Y+EC0Bfk/LzzoYJER3nx5Ya3pVYIFQqfTHsldvxbLpbkovgsRJ
fjsQMWPiw5clIL078LUouIXseW+ldKvHmQENMO4TNGPlYvVDZIQ0Zhg3HdIDAvn4+LOND0JpRogZ
9DbOp7Q1du70gbYTWCocRQa+PQ7EoA0prQzx03HWB6p5I6OwpQHWJt2cpgGqbn0H9aK0sSbp3M6v
U+u329DQJzVakgYGjifQXzJRwJ94AfQ1WDOy47pEh/Tt90DwscJKOOdE4e1yJTiMMBUMubeYg7Fy
AiL1a1YXRCeJ5wqWj2iAny1O9fm/Xk9L4xeY2I+xx+2tjt4LuC6Bt0sSq0o9BMzvKU8gtZpKbxC9
v4N0zMZCqCqJYcUkCCdEP/YY6+1M/RwaJP56y6vDFsQOeIGHwT5oQkiQJFWVJvU8/EADrqZvHs1m
VbIIYSkrrwV42EHmTjlDPIqjPpS/nBkMpBGkTaUpGuZnyCtQ8+xABxuAuKfdb8UWklPOXjxylsnw
HsLXhDl67J2AZvd8XehhTl4RLtSWhndLNCJ+wUQu1RSkz/686kDucokUYJUBZohrGVmF82DT26PM
+/CR80EuC2YEKC+UnStFk8oBJX5KwE3IfxBz2NZ9b8hOFeUqvlz2g7XJrc0BPCjoQ70hL0Xp18CI
gwPCptHIqB4X8dT4qJcvfLFfmlm/LCuTZXdX4nWkBGD9h8qTGjn1tjpDzz9XHfXRi51xaukQffY3
WSuwEsxrhgT28kqLhlm9nRdt3mFwqQVHbBVEcvTyy6HV62sNR92CSE4xsQmBo3T/7Kw98RHO78QI
sHokzMw6ycNhuVZBCqg/xsh7leXaBsPA8qZ2Wp8C6k0pQx4enUB/rHve2U+BM14MNw4lGF/iKr9I
ZwynMQzkA97WvHbCODOmiW0mZADIEU6Rrtm9vygSbbM6l5nfmc0dBJFiixDq+C87XMGbhcQKpobi
kGoKHX5aoHMaj3kMeXrJUIFfycsUgDSAnTmX6C8pIauskdP8541kFdndTNhwgceXwbpeRXJJGKOI
dbeBfmDaUERplS28T/eiakje6nINBFBNkyzqRiPIAeB+nZT0z3z6bXa3t0RNF3L12D0PlM04CXeo
dbsxbCKBDQebgz6VZAn/ApaRr/ls2L0Tc6N8KkfpRyRovqNv1Mxtx6hZilgUVbCRS3chi9JkacS6
sp0jFFMIrcRweJ/1ECVENKNKn/9Qcei6b/EN/D1Ig7aQLMCPh5x0xMW0X6hWoITdD98QdHZaMqb5
sRS+Vp/xrVSPByvbnilTEIFCv2Karie3/BSQi+YLmvtrmk+3V+IiYbl+DL8OzOKfiH4cXFgicvdV
zqCFeNymRgtV12K3C98W5j05Z7ciLCFz7953ugQUaokwCPT9U7hnToLGRNs1bR1fMXwPnCeFbR3I
VFLBxUMsMrU9pzRs7EqQ1CzoJzlO7eOUdfjWAABSLkp66sYlcHlJ031rfakJJIMP83GyOfuypSuM
MInss0SZwXmTAlhYuZpJ0Io2AtDl5VSDtP6S/k8j7zBRWoKtVfhfaXA/pr6MNglLoh+0b+V+jYCK
xUg/ng3awbomz8Wj2f3wgSNy9DEV+9z7ocHaTUR+CIfI9TY2zEAJGK5FrQrkb+N0GBdHIluEFAU8
gZRP7bNlGpDddAGrBDGyk9uLGbTAccLH3n+j818QD5JNzxEf4zwV89EE+F8Jmnv1OQCV9zcFEhCA
5NmF4D7uTYf5/DrdWOxxZV91KPrCPHL5WljcEV9NjuN2/KuO7oXDspzBSRv85ie1jFHjiazUOhia
jvMcFYstYPGYGYg/ONlTMuKtoF1hmuq4m0d1Q0Wa0uuaCZ8F8Y+RBHMUoDo4nC1defrJ2mF5uaqR
mJW5CLrZvu39TTeCfA+EHV8+MDOXKUtwye0/QcT5jEh5IsAswJrMedbts0nwG6K5kpNt9KSGEWdC
qwf6++z2zMcRzjqwa/6ZvYwvqkqbTy2nVXWSA56EpR2+dEd2zlZOfAaYRV3pYsBBUXdJGLeFWiX3
QHRbT2xQxzXaozzYkLR4gAzxg0W+j4qocDT40C/7hYae8XuRzYxWa2SLCNC0d9ra8wWoFMusOZJB
NVrOzelHGFoPdM4wBKQiFNzZKP0u26e/jFMMm4OsnLHZ3GAc8pdNq7U6v4Z35isSnkuJbVkqOcQL
JIVOgc0jypg54avKz5IJ7Z06NtpQlG4e2b0CdCQi2MI+tPd4Jvm+PZntaYuBZk1y6/y+JpTvSWqj
VL5wHSGJlwuzKngZ+SoFsqH9vn08bgKLrC28oHuhCm8uYbY6AGO8KzuFB4J8pB7srsrWDs/Yf/91
pGfoYpQJuMRkOQ1A8E181wjKzwPVAjZm2tATHq+qDpxPJq5drtST0jXibG/ew/kGIiasHV7GjZ4H
lbEOI47S5sgKfeANi5zPvbk4K/4X4eim1DmWazQMmnjEqC12GgWCwg7EF5V7qzc8kHSs/QSHH+CQ
oQJiNkxV554knT1cBh6VqXQIpern0O7EzvPyikm8cV1OnBv9Q2FrsJEjuErO+YVih1oZ7fbr2eMc
Go7X/gHBEaw+oW9O7RN/srx6NnWuP5GBQVjp1bqK4GBFuebWG5/FCy2knulg9/m0UPExEZ7LUEST
kZSU4RohW1jvhINWNZ3rgfshDocviwW/mnFwCId3xVVe8daAlNLfmUU+7pZ431Dfx6u9R9wSDsBS
6Y1qopiq95d8YSgd0u04LR/FQJSwqW5WTARgSuXlCqNCIXF+Amb7ZXu0dJbUsaa1pprLpPgDup8N
8ZglMZa1gg1JwuTSrUXOVcXwUnTe2PN35+GgEgzuRxm2T0fuH5KedMbCfkG+J5D6gUC9ERiSKOwc
q+nPKCncC/cs46+ui5h6dBB+1pD945yTGWznS9tId8XCthg4qoVAjwaeW3Y+wcHUpMBkBv9Y1fZu
IQpCOhlHdt8mFCeIVKATtkl1yLm+hOSQxPuqEOTgHqtjXlchdyLSg2+aF/KsoimrnstZb0oQJ9ak
AGWCXU8b9plmFuvU/R5oIh3fIV8fst37kSeyjGiJ7PayWN86CeH2rqn0TKhH6vi64hkUykzba+yC
l0JZziP//vP0kmQMa9wpnhTeffKZ0KphaEglSVFb5we+nwmBOa1vvAARoBph870ZJwUEfHElsU7Y
xo4PsgSY+ArTiIN7XzJiMyWYHgu/JL0U25ALA6k770WKuG9Vaju99V3NbcJGOiwVpGVqxMBRCuyt
g+qbMZUB4Myxf5uvWYu5VWEYwQnohssNm/1OYQf7BMJ7EqQC4RlGU0Gz4GGXUp2kDmDeY/L519ST
u7XKor0v3RRQQklZjc1WE7fvzbRw1znq7hkgnlQjCbzSDZ3/3M5zwLbz2kru7hDFxkzCefn/QeE2
oiFbudkgEAaYW6uNx+lTS5s6JD2qdGzlNWJSTtE3xbx8eoFeS6dqeNBODM+1Kyn2exy+U1jIAIEz
KYFU/+nRNltTkE1215cWSD6VQJjC6KJJV+Sh12eYW1gUW6yICOGAW11vQZtmpmbAv9teBCsj3oP3
IJqwBu8JcnxvJhvvbFzi7QU8sNnBzQ1r21Ctb3xq9iR9DuH2yNdaNWxqVVEgtKplTtAHJVHKp7an
0HMd3/8f+O37SOoKMrD5xvdlekNyi1x8iG9s+IqmjNC0L1k8y4oPT+3haOzer/0IlCQioHpImRCZ
QPAnIv/9NlLnyIOdZafN9pNgn5B13ROPBnNX3CAcyqFaL+IHWl/pNn0dASLXPCSJg+OhAVmM81c4
1VyKG1U4soBQJcmgUVrC7dBbEO3KZPl8yDsBpKkNgBpxCqKN6wd00LcKETHjGG070bJ5bmNjZy7N
XXn6ZfVvnKBHkNYiEyy9IVL0iTqe52v1QhhrXcZBZl6UIdAmIeRRQyK6zmtJRxI3lEPBqrW/IDP5
tzoNgZYOz8MSAqMA58CfUalRJUDsb4ZEh8aK5eGFDtzDR2oDA5HtjpKWolPp6e502lQlG1rAQ0F2
LAGypuKZ6bv8JzU4UjJ9XCHCenGnmN28uHdxEQZ20FLJJ7IqfaRpm1BI2wN0kOxQFqrFttmqBu7G
ITwKDxzQplo/J4c4bJsuEMZsn2QWXu7kwUWuqxSHKbMmuv6en//9qaU3gPmCIJUTLn2OouRWQCrA
PUjuOoeCEqPAR3Ya2K/6OHYFABujPD6HmdQeRYKvdm8LpFiLm2841U14l2htKolTKz5jonHeY+97
wFpW0936mT4RYmH/pFNQDo6oZGgeUOKGK+oRFyddimqBM9JW1tXx8ly7I6VZ5JdrhQST2fSKjjnu
QhXk471Lvbi3GW/q26zbibNYHxG/eDww0Vv4JnYkgLYvmZ+VGC+3JOkDQSQp11hQo2FTKwkLJmvr
04Gl5nh/EhX/nLC4RUcIoaYV00nKxPhQFV5N8yYWUWRucF3d6T3cgSK2hjr1AoHD8tf5jTC4Eg0I
Q4t+97CcIHZphL1el0l84TBYiRn2ImtpLPFbqZK1gUBMHqlfTyy+Q/aupwWAVxP/I1Gc3uet/3xa
gpXwFvBNhRLxFwfBRZxf6qGRBlPY/g3xrGAHacf1aofQxy4BIFQU2UqrG/8u2Vc4sRe0vLqz5FO3
dAqAvuocXZLdcspKvq7b5PoMGDz5ssA6ApGPhoDQI0RV8CBovp8DPEE1Pcq3BxF8We8+WICnsfgL
JSNzUsETIAcuochT5uY1yn+ooP6OscpJp8hriVaz8ECqalAF0IepZYvXFI+w8v/tHhiNJCvn1axb
BHgKQu611lFYf4qKesDzKgf+PLnyekARtbB8dVSxRWMCz98xs8asZA9Yl+nYIIrEiKGqCkmh0kT8
GMY2iRp+hqOZfqMLLR4vTaazRiaKgmMnbkMwsMi6UYlRyH+6GPsSZ6eITv9nCJ0HI3o2a6kW+4Ja
tIcy0XFStx6vdNvzMuxZOgIcTJVZb2Wjlb8fe2RAIO1THMgrLtgZV+nr7cyoPxzx7oGd9HFivms/
fAya8+AxWp365RWpqF6JrqjoKCl7Li2i02mF8hvbmPB+t4isFUjhyNznxDSr+aWbK3sFtX842oGQ
GeKdMFk/vRZ3JeZd0rzVEDsUzsiLNy1YcGjMuRbMYz688JUX5N2OAuHv7fgCZ4HuGD2sI1fe5db1
2jykQPPeYMt1npY58xl4OwysMeVAX+lDFk+9IORUkop3gQpJUNWlOH2poliDRkMb1TyevISGRWDu
5nvS2iL5OdVJH+bYCcWGCDbww1eeGKoSKhnN1VBj6I3LBKrNQD7m1hb7U0ElQxJRxJGSqMc3Q3rI
VVZZy9WToTEM3t3n88C4w5A3x2LG89X2xT/lRQINoF18bldkYBTCAQ7UeHbvkYXFxFCLfSfYgl5I
9epOwj0e34vuzOG16KfJZov9KULd7Oxnti7pkqu/X4XhEVOv7x2188nuiQDl5PygQuXKkbIqjuEc
c7GePuVf3Piw+yOokQfVSnrDLT98fk1N9FWIBI8VQRB/6mabMWUa1qv7ugFUtI7suxnStQqbylkJ
ubJ27EsdIvbmpqPcXxxzqoXhDdfIBS0gLBAqf2YNEb/2DALOzlarJpIalW3Pph6CB2as56+696u/
KuCRyeORxovTOmDOKtghj4ouAdReyLOZfXEHW0JnSx2TzhNwcjiC+8sHfZS1O7Z5bjXECy6QFADk
xNGZlat3IcRqfD047SSYyDEjlRFerql2ZeHXBTZNeMB62VqCfM3W0mzIOOwkEf1U9xXYbR2jlMOG
jXsS+mdrb9QlEEv7609XlKAtKbh0R+r6QBUI79QA7wFnoUktG8fpVL3kQMPxnqNLmlp9mIRZ/mrT
8Fii5UASBlrX5lM/3sgiji/J6ZXhnAqdiYskUE3U1rlX01PtcWhMZ0Km5fA5al2/gp5+PBmKGT8Y
hd3klwGeAZlr0+NoRS3O8dQh8yBFkKWER5QhghDqkQimXvlMx3zFHBXIH+YPKSy0MKRkRmL3mpXb
r8Mj8+9GR+87Q1dpAifDrZY8KJJYS87AGOx/EcsYTxMXJ9bx3P8b1051QqEFoZZgdgmKPMoupSWO
cGNpERTs1FbLEEQVo9c/D/MczIY4vjj7nzTQCqhGyAcxP4LgczHHZvmL0cqGEv+hGQDFATnLzpLx
0G05mwJzZuKR0jIEbtB+5ZIG7BzpqtFUH1zZXS1/3+wIPjbf+PyTiWIqTDYbTVF1Frflu/86ZRZd
lOjqaehanQLm6cDupCF3k9XZo5/gpBZugoSDf9HGtGOgCZuzCYR3Q+yrAXhPrgTwmUqRRnELyMZm
6FI8iYTU5HKKxmrgAn2O4LmnSqeLt5/+/XCfLcix8dE8SXdColfVqXhhlwPpgIYzKdWY+eTqbmYF
qEoTH+x8Zf9CrxM9XPTszBNwmxWZYROpYAzJuIfs1HAa0qHbbHKRFDvIsnrs1XSAiLQc9SaBRdei
WKnG1M/YULPE9JUxJdDpSjC6Sw++xMc/35eKlga7Y4xLDpKiV+dKPmSvOsIkdZ0men0JcxbniEnK
ezV42+u0bpyvzWrGtqR4pWXzqm4Qurqv3wtKm51s65AC2kTbkyjUPrx8INy3TyVyCEBLLKIr6VSD
HA2VpdCY60CviLjBL8c6TEjXYSLlLvoa1WMNFqSSTq9JkfoC6Je4wOSpEgedmvD0S/peKSOVk4vS
pt0WGzcs7CjKpVqpwxy8VRG1rOUHH18gMGBoDJEDBsuNDnMp6re3e9Tuj75rklGgb0htxg2eZ3Ds
RFyLOzDRowb3Ce/gS7aREagHfqCo8VNTYnt1AOoXBrIkCrolPsxEBKsowEvsJ8VBK29mAqiA+EG5
YLwpFG8HrAsNctnSl478phQsP2oOshtCGMs1ZRcoUDHAGmkOj/zt7npCn12QUu7ZzGWXp0RpCbIe
/c/dgJQm6MaeBmx/rd06dC3WmjDcJ+u+iumjZnrOmylcCRNDWhGeY42nNgXmBGHFGlM4SC4K7eYf
sdOogsiVBErp+/xIvYr2PpaYgpy+gZgDPpnie5CEusHXVVxJoCE7s5z3OmYhbslBSNirtzARGUge
TUDARdmdLeraixMl45RMfWCZUxjbEnG0XyKvGBI9Si4a+SMcImmGKeo0QpT91wsNXCobNqV2X5ti
jJyN7lTLWrKqri1dOYSpFVZ66nnOalf+UMsE638l07XolyRoeUt44RgEYv0MuQE4jj0leW55JLY7
3uWi0YDNO+WS4J9bh/7z0WQwx30Yu4zlVPW3W2uC7PzihDOXTuiqFYAuWH8VFEvIh9F3LdIa4XJ3
vCJDJpvGy8q46VTgC/wxZOdpPAZaD++mxF0pZ8XSzG7e8XM3X67NEoffGVbRTm5GVd6SeVuar7Yw
P2k4+DBbFBTMq3MnM2wuFxfImOetMTIM+9fMhxVVFnKQOReRzTSHxaK2tzNUPY0LJwmk8+DzQ66X
SyQDA5MQqXLaz2vKg24B3z/QGYjj8WgHvBle6tqrsavg8XZy2SzNvb7BwUKULD44O/pqfXXSSiZ5
4ozs64bTajeENzACxpZOsXh53iypTo5cRgkEooh9dPMCGdUD2kkRH3XWglUoLdumG7W7X8F+NY75
OgDz3gDA/gmbchAPrm5ejFRAa/JXoItK1v9KRM5DPmMf/7KTOrmO39VILs1bezrZ7j7tGlEi4hOh
TvawzB9HxNAw7p4JlgIbZzI1kFO2ScswhkyMiq/VPMbm54i7qnmmiCf3hBYsKMFZt8f9DumxRZ5e
37thWtdjNCTi2OMWr7XbMzQUylrP9iJzSyrkJXOsJFEnjXRz6+Q5wK6C3OTVUYnpsFR2JLL3gYAP
MBidageUVRtMvs6KEcc3FEssurX1qMF6C/4/dqFu8wCk/bH1oIjht0OibfKV2d0/vjQT5p3rLkgV
1vP+gD1wdNP0726BbYUqip1xuizdqs/yeED9Dq2etgo86T6XtSzhkKnz4kLMAteBmm9ZpmmII+Jn
fMg17vCMLxMLy8KZ8ZczNEMEzSl7kJuH+VrxBGcLeqA1kpMJrytALymIoaKuMMuvsMgAfO6cqnkI
y1Vpj4kb5FIFH85JCfT1zTEcwJ+peNsGa4kh2rN9HTbCBvl5cTGyWZsQylb38wRExbV6WwhF/fb3
H/LupjrlwrEpmCgeZVxumM277AXsRmKjTPqeUB0gnWlBCHM2sjKKj5qiwlXxCNSRBKbNxAc5BbcX
WhJYv9MeAdWweSYq9UdC678Q0Kl5oviFj9Xyz3QEiP7Pp28iuYio0DrUQgwO4UMdjXVMeIcTepR+
8Q6L66Po7tT1RzWNJlhkM/HKOBFwiEPZmAjJgx01wQuMaua+js2DPBZfyU9cwbo9pNVUMWMqAmWG
xjKe0JloBUnWxtR0f0g/5dzeHyPXurLIfDX6ik/j07EdyzB5mWmiaRIua0E7BJc3vpMxQ1/T+dpG
QArmpqZ+DbQ7bQLqZ/K6CDw+I3Z5aU+rxZ+EXlYtd+P8TeGvs56oj/P0j8iFzlDohHAY+rykAQBS
WQuF0W+g0lPQcuSNxYrJsmESwJ8QxJtaz+diejirRXFSQzjbwvW//Xx/ykf7EhuViXXsIrgkbqnB
l5iE00UpYZm9vWH+i3eGpa1e+o7hW3wBLku7eS987OSP5vwOkIg2DjPxkv5SQ4L3q65yh6yb/IBA
Q0LfSDxzynKYwFYrkdI9a2pknt2Nmg/QiNKu8wftYJNITqAFPvI0NhjgfYMz7yZ7HqFoxB8wozTF
Ibk3pSl+TwiwisFXSqIV7AtA2Y3WQcwPYW3Y5JMBongIPMl0lwL0yBVhI6bTWS2VQFrkGW7pg3Ie
OZiFf300VrwmFb+qxoQjazVkxa8Ptes2QjWNM1TjcqM9MXgoD1/I793gYZODacEBSVE0yC16g2Wx
+NrWMfMrPqXsejBVBGiWWoe5TGDUEaFMHPwGwcR1URUAI/15ud+1CTCvHvX4jJ0Cn2ypJf/Ut3QQ
dxiv1TZ7pUPf2Yyy2Wwf5zZ/C5Z6p9Vz4Pb3zYs3j6aMrOZgaUAjDKY/lHUez5hKzUn7T0WFzDbi
+LxV5Szziv7GGz6dtIZfCTaIEmNDJQ+2HK7qmIULKIryHp+3PXrcqYOTMPBXn92pyKORaqmN2iU1
eY1rqgW1cbkg4M69SDJ5h1Vcz6gVxTCIyGOWBzFsQds9fX4cwv282X8/MgkCu8rK00ihxjfAGX5/
btGq2eOSKmX2U0iz5z8zUczt7JzWBfh9l/Pe6URBkQmPSVH+Nqx16f94MM+xP8OIvzwW2uCtb0Ax
ktzXXeJMnkn0MfSy6ASGRM0aCnVQdYmZ7+4CQA7CcpaymglywKQx2JQVt7OtXO956byHtEyRB+0K
hvs1sti2LvSXb0OMVpKK4xWgL8v1x2asuA8ThOgyzfUdigzhT0kNxSNlr84je+hbSrRpvRazyZAn
UUqTTq1puGX1xB7eJDeiTK9Q4Nn9n4x3yFbsIFQa2t1Ka/sfKYTOfm7NWz1reW2OTPFhOBl86Dpw
yzxVcfmLDy9/CLp4p3asMejjTQK+xAOEyrZ+KC15YE94H92S1gFEkuVXyZcllaQFl8vIT2b9BYd6
qyXPI9Dl+prEj8qWybGWqhG5qZai7UdiU9zVeWsIuuWyydmksQtc88h8LnOzBT9gjDeY6mYfJMMg
oXc4hQIOe1RxMbXPB9tnbGdIcoj/3t7GaBBs3PiHK0FpfyRS8BepQQZ+CEqV8WPLT4p+ULkSs7DQ
PkrqSJQpuDkVsOAm7VLwhw1eshUrymg+tNnNXP+uYy7yd9ykpqyyhjWf3kF+mmMrjMQ2kXs2qLL3
kX3DjyVh1GghQYOU4y744iLH+e8FRV/0s8xj5a718IOpld4tvdcStF0iKk8VoFwb3i6amnQMZhd/
xG3tinWWZRBcAonpExi9DjXlj4c3ekUlBPrK3d0D7htdxO9+kryxxSHgm0eGB+gXFkpjhDRg/1j5
rUWjyupO90VoIYYIBELFOFS/Rx5p3NxovxlxlROHqFAv1ZuwOox80KTjm/MKgb3nO0WpZpYA/mW5
UfaEfgZ7OvX9yJki+O7i5rNGYd9DHAOWk/LPldvkE5k1v8HDx6dxY8ozVyILXZ51jDxd1lQSdtm8
130SGDvnW6U+xd6WZvVxnh19OZ3kVQg3T9ar3f+0qEDX764PB0D6yQ1jBvoPx3OOrL4Ds+mAbtNm
uB0+dIx50wrY/Bn+T7i8nhVF952s+nZz0mWd7PzBlKsMoDG/YdnFtJufy18QP5gKF3htfVpJiYeJ
2QBYS0itZGsCjI7oEgCOXVOGv+niGRuo8xgfym+OnSPwpQ0paB2uqIUge7WA3qcCrhTGr+j9mMqa
7S9UaEC3SE3eX9P/45OQ5zZfqHKNjaJ3lLL+3TgSXSrbGvEZLkOB0O/CO0bTPFYWHKhlDSQZw87y
JCPl+26E58ExAu6/jbbvXq3m4cHDrjpOpElqtU3IRih1Ebv/0MGqgTAAMLuHVE0QjceVYc9LeJg2
UIrlGBm8bVzhcDxsOf4zX9bpH487XumqWQuzJtH1yOCPt6zzp5zP4N3J+rarweKwBZv1vvOmI+eI
2Oqt6BhlkRf5+wqq3JDa5P4ns1kEMAuF5LE4SYuHgoE66ixgkv9YX2EB7jtLRAjhmNve/yyJQcH3
4X4BzYfdTZ+ChNZhL6nb+m+CekCAiCSb3v8e9zzG9qetl8FzsLh79h294TNCOJpeHy5s7NUwzytW
geQLediPwN2GOpXCh4rngK6PwkreuDQdbT3lrvaUgBTHjOXqSCIs+5O118LMMTe/TJO5nurWcbNj
n62n719+2OF2RoimtPAtbnM0IVMFod9mOFoDwxYwdAc4Ve9LdwgWwK6+6qjIWjtmdFhifLHm35RH
mY7WYnhicmiVkBDdSyIqrx+E5rIrvqj8c9Lv5bZF4fkkaqxd8/YzndGPWBy5AnYbrhzAdfmids3x
60RrGoKINO9dlGBwqE/jjO4+Imel/vrAKKcxInzIXhqF+x1MNI2+JyhneFN92R3kJlBHrwKWLBOC
QTaQo6DC11mWg7ChCWF5knxrqEP4jQ39UlXHfRp8MShlnB7w5tAjtiWs3h6lr1CJx65LjkB1QkO4
sMMJ4eAA2FSRSiNtAVzcbb0m30ZsreRrS2C4QxjbXQqNkr9fY4mKcjR4CI+1sfuoigyGD9qISrrS
w2d59gdcPPqy/0FlXQEecLPqPM2qidIB5lS/UJU7qdbzeGzf+4w/9Ecy4NcigD2KIVJSo3QFs/38
6eI4CLGY2ClnOBEJ2svd5UfKHFHxH7pTC2LzUZvV+hd+eiYl6ZsrT5AMFDk0TRTphEUgKuuZQEz3
jvJYeBo2GL1Xecig96iBhHOOCjUXShVR6CbitSXJnfxWo5dAH/JvsqZ/yZu5+LdrNDbjt1ilCb5B
IuM+oJKxpotaPtljsEKfCS6L/LR2BXERASvRTp/EAOH4EXnU4aMWO2/GlfQO4s5uzO4wT/XXo4mr
ecDOGqM4D/1nkvAP9sUeIGhKqEMJN08r2j8he+Kd0b2xBe+B4bmO6+pCjXf9R1uYV9v35Z4cXnkg
LiXoqaLhCqAbfcEz2U6wJAx63hBjRse6roi0U5Lwe9Huvu4D1FTlhRR8jzPu4WP5bjZb7RwNxbW+
mC3jqcKbmgVI9e35RxfWcEq2wqqxoL2iSE9j2HWFAMO1RIOsDVgVEgfU5Yxa9WbzrPef/2DozEDf
c9/FJ66fFzPATty18uhETeouSUoucDyn/wv7Yg06VmVTRb3wWKXwIJt+SVBqFkIJvigTtTk5woif
z+2L8cMv4oeHGBCb6EJHYo0s5dUIdIASFf15jA+fIOwYIpbjnobYJ8ucX5BAGuLU6ubcL/XwSnvT
ecBSwCi9ZYGnNmWOyRc7WAZhG/FoKGqezz7bl9zucRjvmnfhW8lBxp4d1+1ofJZG9CEBBzMkLmXe
BrWzkY4Zb60HO4laYOeRkB0LEV8At7M/YjZgo18TX9YBA/6tJqTjhaW6weA1b2eG9i3o6GKGsqtp
gZXDvcTBcVgfTfyUZqQhQqthOXx6o3TdQpzY0RK07dw2rQYC3AOjpjGe/bBsb+FSgSBtcZelI1+9
vKI4/m2itJ4Ed/g1A1z9LNWMsYurfrEncYR9/obtJND25qGoZIbduWXjEmJ/wIhEuuCTxT6igrYw
n3abaPUR1IYLhwTLl3wPfzGdA337prPMpR8BfseAgaBz0K8PIZdOq58/XgUeCVqwl0TJjI+QuBuC
uv9mrNoZpntKItjm8WGXIDLHufFJaQdKhxUKjkoWwB51kzrDR7ooKIU0vbyL8Z52f5fruwMrHwqo
Y0fU+0Qm+ecNtntvQReN8ZAgFEA2SYUpwaU91t6roAoY5v8Wq01GiZbOeoPDtgc0PvpEQFfzVakU
ee/L+47FRkNoGag9cjSBAY9oYR9jf4f31wna57ZsvvfdKDqHBdtE+fkUIWh6btiJ8tZ/ClrYdN3H
aXrZ4672u0mk/N6ZrBaooJhs6Yjb7mhrzrE80VKWOzjuPJbx4BMSajKlYEd2N+P0Ls6dNGS42S6c
aSPw6XCJWu0YxSqfBYWMQdZ741flvGwkasfIvYPI6KdrMrh8xqIiUdUWCt0T8RCsVyUqrwddMT0B
ErOiYpY5EC1AyS+gmXBFZgjwrCpFi17yVLrwFMLZUwAQ2y++wqf+6d0HRVi1xltvL10YqjHYVELr
E14Vx/IF4ErFUDBqYG9WV3QzRRrwt4Seow8owgKEZ3puX8SDhriY52aIUX3mOKcXr/9T9IIlVn+d
7iDpMZ+q+4/YzOoSjW4k0ym3drpGK2VnC0DJTb4FqbqkTE5QxiiylN8hbnmWdMwkzSnWH8ds50cm
bND9ugDnwlkH+V4IQPsigYI57ocnc1ZuYR/BP2vDdhk2P4HMP0IhUjmpwOET+nb/7XHRiD9dPLCL
ZJCsBhcaFMGx773gwcTEpCd7tfkgkX1y14lOGqTDag+gG/IQ1HtYO/8qaEXHxv7vo8T6xWcb92Cs
KwGEb6rM4BIL/N5gVZz9cyyX88eSRiV/5S0YXukQOVmUJcLJpWmUmUNRl8dDXkQ0zDWLL75jJH82
hqvK1iBAsTYIwoKkNjGn7+SwC5/7MvG2+0vWGeNtgxDH2b94TMdPJUxmrSzgNs9Fovx5ryrcEJPk
oBlb2nXGOmr5rQ2P2ilvKUI0ebjcpATwuPYSK5g3DnNT+aWrU0G9c8QQ0dsFDGVk0/m31OVJnsa/
/+dZyMBBTXIpM2U85HV4IPs/vM+yMZB0mN2eHX4fZYKGvIEWA43c/6Ox6B2qgbHoK+CmSJ4gyT0p
5a88HAkEWHXCFQhcnhki3KGYVFJmrYfKHd9ez4CsUByCD7IxC34fHEZDp3xWst3AfvnkpsRagvpA
8AuZkbi/5F8U8doJg/3Q7whWjPbJRt5mnz/NLJuwPLZ7OztyxSVMvdXqdUyt58C86vzM1jk+9h56
shhWpwZ00RoGUCJcSsEurbLxz0eiN11UKvaLwEQ7l6Dh5Y/Sol5gLdaJkhDWDH/aqDJDo8YgZcSX
TtZ/m5OmQFD3kAbWsKdNHonwNjBI5qgKeZKhajLJDRTlUNtMS5G4F2nWOnIBWOra5SBfw02PUbL2
yPHl/LWqO6gRQuHuituodQoobs1sbFy6s1QmlHy1+NlSl3aifn83OlhT72Zpi5XTHUgUOEogKerS
0yA4LgblTJ4CrCr3Dv+CzsCJrdVltrtw1Zo2LRg/e3+aE4Vm2QhwdLa1KNXBungaoQ51odGO3QZh
BIUYvU10F/u+Fu1F3jaCMYOdDQjfpTXkXUDCenfCTW/l24fUJiwIZAnoY2kmKJZl0Y7RCR2hbjAe
aWdYtCUFbLntVXskPkAObX0vHm4DN5vjoKLOekV1rN6LalYYou/nJYhjx87N6S0R33sOSkk9d+Ia
urdd1b9YNa0q/6xvk5on9wJbfHOmQ6ZvYPJA6aS951s6HDY0P10Mb3xACHIf3qAnrpWfRDZnq6RT
xKMJCIYrAbOCJW46STo/x2EolDTbK1JUE+Xs7erZWyecmkVTS9X40rQpS76poii0JoKTAKcDjQbr
VbBly84Q4OuGq3T92vZWizn6NfJYEki1JvIvKP1kV7ksWY0i2USKhLY8p8R0+nxWcdpeB7EB5hDt
RWddbliYzZ98VGiX9yl1VLRU6Rbl0HXJpv6ey2gtTptY24VeCvcy8l3Qpz9S7BdcrpD9h8jReKUF
jjN3Sbwcz27R998KnJLpGg5MMtFj9TEev1Wthz58DnqapNeIBNAHgYB77fTNw3ypswrljYyoimN5
Uxt1x1eOJ5T4x2lksSvUjJsVfdaVqy7ESn6LrhEZFQDD/VsZZrLKlb/4jPZMfDQOqcYZwt1GCnmD
AY+AiOQVT1x8zsqQlVRyg/9xUrCveZcKSmIWXL4KTH9rLpk8//SRiA5OtAX31T6q0FX8AGP7Ov0c
Igv3D+KbtkyC/BZB8GuvuEocAs8Ch/SjHCKxNDFu80xSAJ96/Uu86LmbW+9yCFNmR4hvWH+eKT6V
b3WIWuxX9LDzPIIrlE8yLL3JyS4li3/K4QnPKJSXWYFlnwiHbeeMbNJPFl3b6fH4ElZkg7hktcMm
lWqED9vft/NacGuFPvY/sTZeS7k2JN4sNzvziY8P66TysxAmFCYn0eamKqYImTLGBS3AnH77d1+j
nIUYeBPVT8RCWwr1zYFu5CZYYi2HfDY0MywDpLlp5249QuvjID9ffQ+fZOl3LGGYaTd7BRcIciw+
OSd2pc4vNfix0HO9iHLXnNs2fGfoum4Su+nbeFEneW+mbfmwmLBzgifkk45mCt4Pe8i6sFekDad/
Kpr73uQ4Ew/DY2O9fBFNCUnJiDMyBG4+azIRCwNOQXrjs6oiECRLV6HQ4PxEXfczWimCr9CN2PNd
oom2q8J0BfI/lEOdfx02f7qpoeerNvGpjrb1DyTIfZqo+ikjVxAUIE/dmEzuncTrQiz67/K4VlNj
FsndXNO60PCxLL1A6mNuoL+950Yp3LKSMFu7Dm+xuXW+9LHiSpRdk+onxW7un0QjEa4modKQ+yAY
pN9Mdm528DE5aCUmWdvJnDHWWY5mOkvdfvieyMB13fULgCjAmzhfwRkNm4oXDYtTv3eUM+ZMBa+t
Jy0PudxvEHbTNCYltHYYVSu+tTdbnXEpI7+mtG7l75nHRTiiuSzjprT8muEST+FySvLnmYpR49A5
tX6m/ArD5kfxBJW6nIOyLUO3KwiWBP8kv/RiGaKXbP7RT5JP/NXnZTNiE/0szDDVXsNSmqsU2Sau
BYiX3bpiLVmN+jj58lwBsHVKFBMuDY03yM32scf8wzl8eeHe+1f8sNV2M3Jg55NSY4lgXLAvjB9Q
cNAEiCxnrOlzcGh6WkyBEWcvVd+L5m96aO+f9GM/yl2f6zf3fxY8E0//oFpTbNcX2zkVICCoslb+
0y5CwM6BAtbl9rFHJgcErgRUQCEprhGxjF387q/k7nSj6MrRCDEy2/R4ai5f4tbwE/c9NkGBKBrg
tDOGh3wfMaZZZvNYPBb/CRUP5nci4Lh+93PFLKfPzbK6E9BwAqrfVY42tPkK3804+2v9NX75JYJj
M5U4I1QXmtErGbLqUgPPHwPosKSO3YKL+GOYYVVJ8qH6CR9uXoqjcXAah2cNut3Uxaisccss2Ttf
bDdQ/AafVi0Csw0Pgd7hVaN1g2hp74isaU/gmBzh9tAH5faQhwJk2ZlxZNIgDIMYUNyKN8BYNgoA
uxUMAsiRb+GYzyAduHtZMjHsqBV4ENxGRb8gjTCjiGJTFt2BenHhzSpQKGOSyQ9dDUAnKgxAFdmB
J5m3v9obGVBpV4GE2l3fyxFSaeMQvDVVzAiy78NnQg8TgSzaDDFLPSREH3MwCTHruOVxrvfVWkdq
0kS34n8NuTpuCtSpslo8VoqOtE1kVwSBdVC0pUcfWXgmnZZnbRqWq3WeooJ4MwHt638kxfsVymf3
oPTOn7vvkh///91xFxKVNV3LL95INsVciVztn3YcI80xlD5PBELJMT6okuhxsGxC7jX3ldO6NpTk
PKHg+AN4nXyGCtXpy5J5arpIvOF0UFyNvYDoiCcpPYEr4U5heEEUYPHfVLSUhrnlyNyd6d48eiwf
96rgzPxvFw7T1qqklxnPZlpUVvWqz/T9Gp5r9SLp7mZKmUCuq+fzkniaEZp1epHbWnBxUIZ1YF0+
+PodbhdEIjEqAojj31lA4r45aJw+bop7wpr82Lnm9BQag0qTm8McEf77MDKLsHxpj5eVICQ7hpqb
eainrXsQv+OEcUKGWTsu5sqVZQKkyv5Y3zyEQ2SklQWHM2+NiRR0qam4JqWnH/mo3+aQYT7PlK/V
EDrj/w34giqnR5L0y2WwsUCpgB4F4GCOXZTndsRDtcZapNjkFTdG+hRdLvK7w6uSU97rUr3I79Vu
YyM8ClJWv79qAMEHFXWQ94tNGIAV9y+MaWhOuZdqafSRAsJ6rp1qFqGg8QYcvQEufSLvLRw99KhY
1qJA77BwIOek0VVtpDPabn7GkYnsme7MMi9cM9sRfoErf5HvHgxAGaHx5n+IA+bInhZ1fRCOjIDc
7+tMyJLgueWlDg5PHVHnv7GRinziSGM8KLv78uKnhZijEQUC6liTZZyHiEoyM4Mc4JxuzMxBKd6W
U6HpdMdlQECOyBSj7Hb2N+MqSwEwqgH//SFqbWJ34h2HuhDOyw5Vtkov5IRO5u11OcVu2H2sC/Lu
enbRZr81BOhrqzAHqhGaPpANBg9cgwbbkazzE2BdKzfOZ/sLFJZDKbjUBVperlW7fdI6RV58CGpY
1a1u9D/5xeRHdUnJHdqBRO5F40zjlZiiM85GHVwjjJ/VFaH8cCNSSU3YWJP4yrS+1rEOXY35MuKA
M66nxwi1GuEeTjf5w0YCPfDg4+sJTFkNDtSLOowaT8LCiDe7cjWI4trP0RdlvRHFWCih0yH3F8Ym
6F5CLn8uweZOwCoz2OLdRr49EY/G7KrtJiWq0fynCCFf/fJcV/UtWyrbwIlxp+orRamN/fdLhhRR
mpuMqQm0D5Ps+r6upXNkVg/KUfxLO6hg5Mg9P6qObaqCBm36u2YljBFPcFa4weY7Bh14b8PN3VDe
+Tsk8ZExORJDkx8jmwlJ0rsNacEyz/ZyFjX9c3lW0Ntv0XmyLd3ChUaCaiHnLK65NS6R5g5BvFSU
aQRO7iApVAN1HBA7yDaGCdhT73mtmK5D9U+HMN6M6YeM7WnXcF+0rTzOIXMyOwzQkPWCAatnonRS
Q38h9J1N7BtHEkMju8Kem59/PS8ustB37fmqsSAfglCkXywHXKyhVoNaiPCfaRlmDjVN9sUvDa9U
p3lOZGB8ZQ/F0D5KyxN1g1fsN6a6CdJAUtlgXl6j5kv19NQ0YXeSfnqV7spo8xQKTS/TmRMwn72h
aGgqdv+wwLaWBcz4royAOp4xmoZyPukRsqYOdkRzci01ikMNKbkk2mq8I6etmCxSHAxoaXQpo+7F
L4b7wseFiXfUoUmh0SbZLsP7BT2xtJ9CjtLB3Rb5DiQu78NbCex1wjd2zx03bb3XzkXO2oXeE62a
EJdku9zD3cD2uZpaWxiipk9WSIka25qf0NRl2XxJUTZWcv1JHpFv4xpZ6++mKbvJWl0wiOjnT+WE
18JZDhhfFbpkAiexOcNPWae/S9weN4wC22GAk32mLlcl7ufxrw5PwZJl5r/xFeSYFYbbPR6JnATk
cAQK86dRidAWp25N5pbAPjySfVYNHBgJyqq0GxXzxD+WxE4z+csyiI/MSIqw6OALWJXjeiVY1d9I
wLbX0iw5nZT4wPm/kPtf6FA2/dMOqmjGGOGPe5K8AYq7L1MRk2I3/1oItWKhmZpsg+KaOLXCM6BG
28QjqvyphC8Cr4q2zWShroN3ruyLf4AMAjgXktMxrk3pWRbTyS79cdSahgsY7pw/RzDsKSKmU2ou
sS0tbtDQOOk6zMe4QOiJt7PtUiWxURk7zibW7yX4y8QOygMfyqc1irFEiuilhoOVcFVZhKzBtf7f
r7Wf9Jx/JbB+RHQNplrQ7SsMNazCUYXnakXsH2m4TDip+JK3bMhvmrB5UZ8SA04+kfKSWCbqmvVo
GF9bSX0mZOBT+LFzxxA2BzT03fcAuM7z/4u6t2M5MZYPsiwweroUl6mRUHhONIJgI37CfF3Naz68
lXlPHmbJqWFKGCr4KFbiqnFqb6b68iw0aOU1vgmRJ8LV4hKEGOqjKgJcYRYqFX4xbxZnABzb1aDT
HAUk9sO+aoMPX0OokEiT41tSXuvnyBZ/kcJI72awNYVR7Y0TR6J6y0YlEIJlV8RuudBAIiz9mbNF
HOODPF48ZvOv+0B7ZoqiYA5ue5WYJmgIVTgywnmE0U/tG9LXxGzhdQ57DQ2jkLbvlbh11Dj7CQQX
uc/SQb3WoXFWXjCXVGbtAnqRrUG7N96YFdnsnK72i/hmMZsCJmFCQLs1vZVbACH++1WGJTVAAX8m
PXIxU2XtH5k/+9F+UpTkV55GabtVkELknYT/BgLu2PDkpuQwgGUuvdgWYPcG9h64Q8pQAiPtPhTj
uR76Jws6NYhjEmsH8Vge9WVXinsdRnEOxZJRNuAk0xVnuIb6evurXMt/EHuSPKpTDJxeIYycympz
5cTB1FrR3PmYWVhVCxUGZKoJXgN9/N6XM1AnD0eHy7VclM98phX/gQ1NCumh8DffeV2W27t4ElfU
lxiJnVCnnWYZFED47PKeel7ZRX/eOUind2HYeuuCrCegt8dmN+cZ95JjDduSROEgu+i08t0RJUan
x3mLj1hCKOCT4hDxO5oyBkNNIKxOw28Z4M3WT6JFobI2kIIRY8KioBCWzcs2cO7riAbB4zNsUgJA
heNsWceykrmIU8B1BW7cTnm7DdUCseburHlcHgRQ4vdCpufjh9tcOtBvJe1A2eJWJYEm86FSjZot
73uWy9M24OxzcLixqIyna5uzYxn/2Zj0FSLiL4TmX0eBLvY5+FmeqTbYgsuMJ/37hZ9zbssdvgge
JHfNrLf4H/9JVNYrbj404W1JwRZRdHHtLuF/NpZ4xomB769KglLGCvyvK4hR/ZXFKmLF+aCHD7WC
jwPf14+3Vark9qVLxMx1IAFpxXbXSlhEPES20d5LMpIQog5E+j9vZfguet6WcPs9qZB8jBSF1y8E
9ievMQJ5BEecR1nvz0zcpOi1Db+Z3FhHaUZnkFYl4JRPktWTjNgZC/ikUwRd/4ZPJZsaDGWq1iX5
/QJTAkGrb7NMO/ZeiMvQdk30GoUw+YPYNfC+CIPNdpq/qnMYOs85J6dy0NGUzAgjrk4MkmnO8xpJ
BL2pi4hLTfciRT8vP05K8pBTjNWDHEhI9r1VW2uGgNCdyT59kA2zGygB5y06jI9imdM48dqeYM3B
jSMPkWfEOgyGEdzeaqsRPdFoGrOsxgj6w+xaZNoNuX/FoTQGMFNluodA29hMzJJelxvhUmXKCSLH
lEQuABfrgsnc+jMI1DimZ1BA0SsRNr9THXrzsNrlxQbmBkIOgeSpelpYmdKU5Q3wPhXUdIVNmN49
D+1ckQLte7N3SuqiDzZnAbh7ysc+HD4YOCLj/lG40Kkza9V0J5atW+oqFf8uzLbbZGicmvU5wOeT
YpfpBZXc1CEGn207q7FZJjsoSkylGWO0Wub2rxPZf+UAFoIE+jFFEyZyJ2OpAAc3Zu3wwstRqO2F
JBVZBvftmVUXh+3nkKn4KBXv7qZ5xSkkTkzJEpKIHrzSoZPZGecBS4mYsEJ8o2k/xPf37a7Y3jLZ
GXV4pI59LtHIT6iYOlIT4Qmp0gdexvImT2gqVqxc8odjP7lZUKiKIO2XKTca5591/McBhkfzyoep
imZ3rA3hZN7gb30EluNmW7mfhjWWheZFg0gnOQ9BVKmgBpv6A8u2VUmFpxZ5qtfa6Bdcp055qz+G
/i+pO9Pkzq99VE8lHF8Ik0fXOIC4r2ga7u/ewOBGQ4unE9sw9OZHqtsGTRDODiraWhakcHfCgUiW
9eaABHyytB0tcMazTTV6PeCL01S7RJp71UsboYq55kq0K5XFqNkIdgj9ngnoCVJZJQlrJYlqbiFk
zuieiswhgVGlIRlIbK34MxSrqaK4G5p48zbvqf8CuiEJdwbpRB1dODpFOoMhFI/rfNqHJOiT7jXb
AWLcrNkD43o6HvypQzefNAifsrtGnxOq1Fo6Ksi8dmrvBsNSX1YBNG0WuJx7Fdt67PqGpBEp+mys
9+PkcHZ23W9AHDmgrlf2Ws7Jq9k11O6WgNo6q7BVKHaQ5i58LnTrns/NoAD5m3rl2J+nokREf2wB
7tGTp7UDCDfcETf7vacyTaLodYG733ZCpeM4jURWBCqJTclMZFNUi2gBERUTjOdV9VQAsUyw8Yzv
280FtsyYfKNrQRPePdb6sHUjmhIEqFga1JZJdYdxuGRoFjQYYv8B+GBfaHf1jVnboujmRE83yqt5
vAOJWTRemgaScKusMlzxCi1t9M9MOy8dNG+ZFUJ8i73XNhtUwJFv6VZRi7AjVem43R/bxgcIWvR/
gn0oW5Yn/8MZ0V/u06pXRsR6i2g+/67NKV5wSvyziB2FEZzDKsghIwcIjOkj1nlpmLbuKsWYdw+s
Tk/1bG/LzVufkhs6nxGVTUTTg7Inq21krjytYAW+N2O89c/krb6h2cNbq0aeQDBzm3VK/IW2NyXm
pDtdEFg2BRVbZXpvCyJC20+yzVLIH6mc1v+tFZEENM5b3gBg3+rK9VRkmW9DcQXk29BeE5aHqRc6
BNh7akL4ijHCZzzh45DTCj42hQB6KcV3l5y9yDUjV4/dBeskXeu2cUmGsWBkw6Svn9X0xTYzjNn9
vNdsgtNGOep0/upAvowrX6x4VRZ5sn2PW8U7TN/fY6bo5QRt0N5OH68CeWNEqqdKGwwmUB1G/E9F
ZnOiOTlBbLc7LUESynR8W8IRoll6bMpfTghPR3kqYxtqMq6TS2NIQBJOh2Xv0tJ7MKtGP+QM8Sbd
VO2tqEn1R15TGUnPEpH1OCDMER+9UThhR4wAC8vC+pKkyQ9HG/omdZeOBimDKrHWCRMYF2B8P/nY
GnCd+LZkxt2SbyuniwAtjflynkgfAi6W/sNeJQyBVbF0fMnFnj99peUH9QvgcoeC24KHxoPKmKM7
2291OXFs8ny3QcGkWM9ELLUUMzEN/Gexkm76SwJLb6+0oBvzmPOOCsg9xxsJyPn/l9pWl6CY33Zg
fB2soC2SiY2LJJ+CnpYoRr9fiv9Of2AL8mYUHOw6QN2FS492Ey//fTVp9pC4St1F6djbLo/mCJja
0nZ5HZBaibb+gN6gDvjrCINA0/mCX87Ji1zM8FpN4mec9eu40hPLiEN6RpFfOkrbj3f1YRgVUY0R
xQRaEaNEoG6gJVTKqPz9hNbRplpnVHyqfHMBkjvWHpSKXAQ6s03/SZE5R+VnYFV5D6Qknfd25tw1
tjcyX/XBAJnJY9M1xY4giB366u+osHl8ZJYOvvQhKmE2W0ruU2EqUUZZn6Ut/Kz8UeMl1P7UbmHt
n1U/RDmJgx8XDMWkYtOQ1J5CAudicscDNHH7DxLGgL3MYTds676ndmvVZxaTq3bRuyKgpFzRhGdv
AtHG5yShwjkE9Y9TEjDkrlnoPEScEBar3WcL1n3W269zF8eTZgLH721U1FFvLR/8R2SVzNlUhR4t
sXpDhggjwDV1wfmuK5BC1vRM5OrD+PmOru6YKtydiJZA4gwDwHVTiT1BfhVyJdstfqGMvuQZZ/1i
Vy05xmp+xsETQ54bfswrDjwTD5TmaJvrNxjfAyonENiWKcjwkl7au4cAXxaLcjAmTAKU/BjNu8z6
ov00ygRRYB0WVUwIwTvkEmX85JrkqIgFk0YSav7dwosKdqEBuVnyWK5/TuMkFX7Qj5TNOLHPivrP
awW4MAD56N6hHGD1uz8BL5k4nuR71Xo5/wsYAQOQWxtQSgcp7JMuWrV8s1Pp2mzClCahLmFOuxV+
TvIUsQJX1ZgbPPWrz/F1WhhZxfe2fqjb8P4OtIdAAD9T6sZ1AArht7CEuzecPu7Sq37cHlo0XIbe
mqucHFPQ/p0FLk+mw1wHL/31ImuVKy9SkUC7fZilHpFx9n4lbHso8sn6TDuC8fHsU81cX4Oo6eTF
FZWDBfxXfJrvAvtlcj+JATblsmAY6YGdrZGzZ0Ybk7UPL3IIrS9LjY8bRR396WyNLxATLN6wMiHP
RNcdgvTSmmW4y+xKg2l9SMEcaQx6BPsFAy1fbDvjC4S3P5UPJWM2C2Hrbl7qVYgzCqoCzEsQ4VmG
MQDz1bE11dUpDS76H6RIE4hmVAq+dfUPc676gRyW+4rS0kAhhT2anZHgzWMKms7aaZpHXarjK9td
87jvFhACVV7V55WkhIEzjOYpUJuy5Ov/YWy9I4XOD8KaJLDV+ji3JVJZRd+MDo0lIUghfKfT01Ep
CAEGDZUr+IwuqtEdSYDrA8PicU4n6/LhN9Od7ZjJdEMr+0JkXbbEwjIkAEtyj9tBt/lFa7pq21Qu
7pXaI8Dexwz246PLV7UaoK+lXO4BhYl5hBZMaxhntzNaIjWfxPwfzEL46e6PtVsVnCNan+TzC5qj
FGyVbdy/7PQDTU9HAkDFw+HDwQnjIFgr01aywf3aELdLZIG8S506J74gNE5gVjAyZ/laGdJxAcsH
sDKYMV7QFAIRoTor2fBDNxCq3seDdpsjK5rsF7qz1NMvdyzE3s//2fRXf0l2znyf1/2zJnNSAwTJ
qXatmUsxcFcCU7DWwXLl8z2z78jsFQbxBC4wriw8DUU/WVBDoSB2sOM5aHlfKUp6XT79G0DnEBWe
zNkoKQjHSdh5BBzZSVLDSWqUmSRx98+jBN/inrZp7wnenNOWK1mTXueNGhExJwT0cCSYg51QQrfA
aiA78yS0KOAauVZX6dOZ0FdeahtkajlWtt9TidzMYH0rGQs+JS00s3USLuzen5iOAphDgrZ69g7n
tWCLma7ex3D4G0FL9jY98gm8eFzBZHVDNKPp97/2JxpldVWqUmAUQJ5xGEfnRkMUmiMAOvh/Lzog
jy7ggU4x3AMIwG6NR3qe4drioTrilbc+/wNXsic7hMtj4H3McndQuN4EfFkEeICe3jwCcgR/Q4Et
nwTJJkGE1BOT+aZzwBKNTR7AC+DSaEXJ0YodplS4C4sCPCESZzIzEKnW4j5UgKx79nsl4TtfLaMd
EMDdUumqPWxbQMN27y9xxFVvtr4lNsNVOfCRKgEH7ZdnCJYFG1Gy8FeyFq0dhuLSmD/swi8SZl10
MuvLWGFZlODt+yGGPMgZ/TCNLse2k3Ybkr+pkTEkSFOWHp89kFUGhxySaWsvDdmdom9qsiszNftn
hsMxM93VtmKrPT5m2QkW3I93/Smg6PbnGkvdT/FT7Yx/am8iydz6X4Js0pU7XI6DAO68cdG/Ak2T
1T2HhCViuyx/wE1sglF53SncG5g/FwOPTvDqANTOILgaj47cjA2bHmIE05y4JFDRPn+yFp+SRJbE
j/5ODssb5hnuw5jO3yLLi/drSVbFxGd17F9uJ0vDyOfQFbzpuOY5awzr7mZ++PYNWAdaoDM5aDku
Qz+2h9KZqZIFctXyGJjrN0Q0yT0v6QSebPnemmH3+ojZHi1wZvwhvl2pgVq27KgQbnOhtDO5xRMP
+I0QndGbmzVUioeJwDN0j3d5YVI0O72jiUtXML1zYkbOYLmMgov2PekgRm0TflRx215bK4WBVmt+
+N93PxB3oczUuP3fRVOwOR14uqkK9ofhv6pr+Uhvipb0Qh8k/tSZNh0i5B2MpR5ABXA6M3VICFgF
fqj376a2HXOP4k+Ydz4lS2cWRTcg0SNw1UtLPAIO8k0wLQtEjjQgUuCAMoy97YHMD68rbEZModpU
Yw2rBn0Kyt8vRtkZ/FTR9Qxo03b1wYg4Dnwdq4LSQphPMGdnoEvk0CFtzPKVCOQVHJFiywVqFyzM
b6ZhuoC3EDYCQJa+uUf18ONZRgvihB2KYoA5VxlbxCsaj5x26AfqQKyfvFK2siKyGAcWkLRcDcKy
jombun691dR1yXR65M3ykDNMdl5nf/JrfNKQnInHz+6eOBcdyWaH5PCkiIFf3w2Ac1OtJawe64IH
NJZpgOxB+n4VfMNPLWKy3sPczi4C/cEddorEoFoKHj2cLdycTVU1ZIfLm5sSjJXg/wuyqXLKzvAr
Tdvt7w4RYTZQF0ijOOP4Y2OmO39GpHqbwQ4Ik5xqAWgZQ2SOCODT6+G7QJ9J4YdBqt3Tfye5KYP9
6GRP4KqggW9TV/K0cHzQFgUSlCoW4MB6oQSkpjNWbqTmtP8b8ivF9DcGK6oJhJGMSYNCZ/Z/ExOk
MqIdfyYqSv8m3m5l3KXRqZI/lLFuXvEo7N0iaN1Qi4go2f0hadZuuWClDCPMh5SKW5ETGvZfYB2t
gR+gHKAGQQ73LspZvvA6ifRcGo/sRTuGWeCb7nBqXtPku7kFQmOol8UJDeAryl/l87f+jj1DZnsw
1qPCVQ3t4uGjmdIEnF+hL2zfeUjnxt5h+18BJoj9uOQC/XH/8MkuoLZfj9dOhWdB0SWay45uGJNI
DYA9CD704PCUvjaGIk7i6gknVlKak/rQGc6E/KOl7+vXTUJjK9lNJ+7s2lww4nzNXye3/aCpOVkp
08/w4yFt3CrRotxmUJy+v+ZgIflagGTL4FNZGNpF7joHRzjKWASF5PtLduNgpqcMFr0Oa0x+s+RG
UAKKLhdwJUmNoRQBEQjVg2Bh/TqW7fDatd+zALbtKRUY1WBjxEPKyA/0jvEJ3q1+b0J/s19wcWgj
M9yFloVpL1D1aUGbJzaRdEZHJ7/DDfY+N44Pyo3PAbL1DY+UT6rylKLn5zB9exPiViMxKgK0dLqZ
RLTARMYRxjLYUleP0D+8rZgL3PPawEJTyjZMHT1AFC4V3edS3Q/wjBXmmUk2cHbrUbBDSf0AVdOq
+evswNkrTFNqyYcZxDhVlWP35AQYqm1IcBaCagDrgVVW+hl+Tms12MNAVpchcVS3Enbzmg/6FePg
j4HKyyepe8awDbGRFp6tl7NeNxR1umTD0fV1u2Nr3NhKqmX4MsH88U3SnsqrTpRDNUMD5rBH+3yd
6cnsOT113i7ZZiWuyRfQTdUHe5dCw0BfKSz6+/8+sFM+rqumUthcfYQSebJ0a32dd1cLNmHEY3Pk
bq/evdn7+7jrzaGhgQRI2Npa1XIlF6z6VRmKbaXmCSDww59KPorb0d1tWwFLwlldPK7CeAPfTTHj
WelIgRCrYBSmLUIfwNaGJsrKLsgLmO6i6wUmaM5VFRYyYfov5BqGWLz7snT9c4XToC1kP0mOgnNO
aQHg4Xu6jP2D19l2S4a18YD35GANvrJvvaGcwzOQx+jUJCigA40DdaEiuneMllP9te9liyNkUgL8
0/kaYPX3k3zJGaOKhJiYyPxvpBWP+f69Xc11wBlbxTuZgVgNsKO1Go4ySf6Ilpt2MG69r+MeksTq
HECSX61dcJ0/5/RxooEKnJMW2foSC5jvifBeSjiIow48tP+VZbNJXmVcqw+L2/1F1tAR6wP4LO/X
h9YwWJzrpT2DX5MngcObk9YfyhD7XTbebFxBdm/rt6uyLUwlUPgZASguqiHp4IsQFO4wI7eTG1ke
OJETpJoqEPULYZFGluDImtjUuQRX+5uF6UnwErEcBqNGenyDOCpR7b3mWV6isDSPA2hq151yK5gs
P1zjbJGbfRofozpEOVv3uvvEbedKbqL8G7qnpDqJi6v2q45Xou954NvdpfxApgypM3YULJvHXQfA
v6pnCf22pRWjjweY9rtlm5lk88FKEwCS6BZvdfYpRFIukjwJJk4bPcJ9auEKUI3bMA4f7Q6qIdTf
AInNTrLpW0TSk9KfqlvGB+QcRuhKNvzyCMzeAFljXvZZ1WYK1FsaOBkGWTcvyaAD/1K1bSYobPZX
0Akqa9nGg02A4bDmoO7MjtzfTkht7DMMyrzGNRViOtpboCSYxPzu3KV0RDGGWdXOhltgKO3Q3DAo
vDb/eMvI/ZAB5gAOvB3dokvySXNQFwl8RTiW3r8m3+RDdUP0j92Fap0KIvWHOw2gDo/klObHzVUS
dbeo6A6Sa4bmBYy0+Mg/smBifmtJUM4NtpvszfRwEZSXPTfHU0mvwtLrANykejTPFlyPnA6EpDnt
LX2nGhkcBkOc3wWAzcJWZBEx4r6j7uULSO+Fv4HviJlc9itRf4niVw4pDREYJqJh5GqBKBwypKCa
y4SUb/SnLJNAxBswaCWbL6vgInWjBeXrbvXO0kycReDLXsHr+Kiz8VHzrt5rtBI9ez0U8PQdjtl0
xwlrnXh4YLQomugYuc59SE/YRJrvVASjO7EAet7G9pp7xHOcEQ15vvAgLXWhTivxnWf67uEkZd29
iU71RuRsOIwqcqVd6ZFEQV7iaaYx5Rw7nLJVexsfv0f3ZxzLhOajf2yKW035OMWo3OYAG96lrkXg
AhI/LIXGHSaAkCy2+Skbg3bntoqOjmqBjkbMhl12Nud1YzsSsN/FlR5x/t7NzB893kvCksLTI1xw
TTcMO4fNNmqSaPePhKAoj6/jXqgRVw5Tbbh7GYwewRmMo8RiPUOC/jW76D5mkge3qoPheKVHWKlS
GGVgSStyNFs5GYg+8JMbneltDJNBkCfNGX6CQ8SDfLjZPFDbGunNp6M6oKq48Q4dyrGcqoRCu5xb
e9pv5NcKz6SaHWNxVpd/8LQq5ZOemWS3zBImD4wKHCAZVj0QgJFiQUccJYKfQwvPNz7UxZbMtpWR
ctRBPFx2tXnYQ1kFie26yu7EoWQI6lzHkbfBfQDTnZIyhcNkcc4p0roxX9UyBKpwWzF+RhYu5cYi
q99GU8zplK3F52Vm4SZYeSmF6Sm85j0NQI1zZSDSPISfa8a3mxAPJ0QH8bSCf16+2/Xzige5B7DF
Y+TP/JrlQxBLWgMQncK2Sp9bMyjAWWdG9Bv4NuGuKth3CQDAeRGV51K5nx86UyeO0rDEB3lXAoy2
hX5ydYzGljMLWFLuW0WJRqv4WRnM/rruoJCKwOTFi8Jv6YmLPyx9fsTvYGM1QNhZhXyvLKS7034q
Ho59t9BLWtEKOXbDr2+ATZdDXVO/VwDICzrlLWuHLb3gS6pj32MwBrHYNOUHyJJXZkzc1w6oPSMx
bbB48isI7B/AizbDI2YbDGuDrtmRCip6GwkKoK2MrCrJMg5Zgcz5vS3YGjOYh42d+whuNuhBL2pQ
SU+mU6gNYydWm7vAPd8FeEgDxe1ZQ1JnpZBnKCH7QZhsjQWvVKrC1jVPALtoZ7K0H80Jf7O8Y6Fa
JbgTtgaU20rVM1vFNnUby+Eq32d7c43H4DSW9FM6vZ923afkn7O+VaTwySXOUf+Xfb/OfMgwkw/Q
sHTU5KimLIAuMFZMjZQBkbQhlvDDD61Qi3BcJy0wrOBstED0g6hotTOEX5aP5TBQKDvCMwWsvby3
jXZARnLMwF06Jt3sdKHdmmdbqNn4SRJ+BNI+39wrEKf+YMyqg01uWdYucW2Jd+tS02UgqGJPHVpS
RGqpBsDIKDQr62pWpPIT5Yu3Xn5WVmEzkQX37BHjGrJhsWxXG8zQ/pQBDRHq85Go4iWS+flK1SFj
D5TBUvkAqSush+zROh6tdRGaErRJHvbeZ46GZrvYZXWrh4YA4mIlM/WQ6lEm9gQT6LbYbUYcy7dd
v7Oo2iKfqHjMMueX7siVPxIOlX7n3mkILasYnPW0S9qeGd225LQJb03D9Ktofbmk9i85/yG8UsVM
4KTQw2xkqhj2qpQk7W1YY/WiV2fVIB6EQRWR69zfAFM0SgonzdBK1T7AMv4dJBr6k+DJKxJ5Z8vJ
Yvi1Od0JLk5rPtp0eX2czd/tG0spLoBeTsLMGS+C44bgnwicKNa3w2o4A0105fBZoL2xJMZsXkVb
14bFJ4wRJjqpgbjSn/taVlVu2a4scnMWzNXUA8Pt0KLY1kKdDd0L3mPdUZAK0U2kNEJDIbGCyxJC
le270dIEGXORHduRqTP2XGBK4v3WXFpIVJW5o7nUnYTUSq+StFnTj42MsWgucYKfs2PTTvD8drtT
znvFDYV240uAnaI64xLQ2rBVdhi1CBtCmJJEauXIBsWjMMS0HnF0HNxUfDpSipqT1xBSQDrr5eTa
IwGFYJjrD+pe6vOV418Tr7pre1VdWJZ0nxJCb8vukBmv+5JeAX3yrGCCwcNAlyeSZc/Chrd/kwEk
zJ6tMhKzWzWEEmDfJTNgRwwzuxY5IHwXvcGjTy0OkLE2iydxPi4RcKW27SHQCkn/2Ns8YDL2Xl0v
zzwFEGDkOrZqlD6yczNeRu1/3kic9QuMkAaMK7+Y2mkv116QChf4gTM/BsqbRFwBHssVS1xezOxz
S9HlYcnR0mMQyIiWmJrPqYw5DCrbxLbfcIdfrQgdoY4/g8FEUltfCzQFwQ0yz41YsoMRZrU2V5wB
cJ0PIKm4SXF1EK2DeAxEi2VULJO5eW5ff1v3uaFQ6zQFMH9bJ6NZ65M5ntZanmvyCb4br6mSrchR
RNiYjk/jTT+lLtbDFQMZxt/7lGr5kDKgqmv71TjXKDV2HNbPO/LlCOF9pLPnajIYPVhf2hzN/aH+
NUXOMfC3/Na7in2UEyRoJU/H22tvd3bf5jewls2ouXiZE8nodU4gS009Y1jsD6AZua1ntVFDeLA2
BjCGvb4q+OSRXejv7hsKJ41oVqb5EAauWg8+CK/LStTGvjXxzYLeVxrrntAHxh1JF7UFR0CoVvl2
7UV1mR4NJAsQu/u0VQR4WM5oP83OlkWBp+5wnWl/zBWsSqoI/danVf3aZTKgketuAOr+evyaZJjJ
Al92pgeidjpmJA9W37TVz6JS/6kSMzzxA4rmhmNQS/qObUWD3uFYtFQZQO1NbelFERZz4HFHMIGt
PvooP9PSS1nsUcGxIPUI7YL8S2YcLjfUJS4z0OcEoi9LXny3C8gbj7NIS55eXpX1R1JTFj4R5Hrq
AIMtAB4+84UXdsGtJwlj7uYF4T26A5UWNXk9wVpGtrD+V7ob/IN/rq5JwNz0ejPbRtDlN9nFVgeE
bXhoMsnapQr1aXRXzuiCS5mJ1+rRpZqM8Onoo/CrWLfWX0sUGyEs1oxZ3aSTvZpqMOgbUFaKGu+U
wQwfEULnKIEaF8bapUBZcU06o5MYc08ivkXWOiHzWKHawIIqMGCYCpkkGKrGmK9FCjjme8/cmr39
HqH5LR6kXgF4Fbv8MQ0Bl1c+A8C6T6a1FcdqQ/4LVEtiAeTZucESz/4XBq3zW5paRu2z5Z6CxfOO
3CiXDMUyAxP8FqLXWx8SpNysuMqiDqFpNlrMVSLgyDabrIDWD3LtRRY5Q7VsKglNIYxr6uH3GuGY
4SuL/8CCTieDSbABt340VGFGycu+1SayNmv/I9SVA0oCmEJLQPWs76r0Rn1kDML/bLahQCP+88TC
5fVd6a0vt4NGP+Ln0QITlAHaf6HMU9wEDs+rx0z4SHLpsbHXMrS6E7tuoUUprGg4kMEWh5M+yqfk
I1SXxbhHyxEVNZlCIia5DmMQP321AO3Y4Imc1BuesHwr48VS6daAJMF4mbld/IGF8sCdpXya5dpX
84sq+UFGNhE8BAiWp6hNrghqMx3IvpD1SAmc5ZKWWNYXC8jppSPy/DS2NRAUIkiqIDaSEFxCQoDp
X8J3WYqj/62iVcxdZ0Uw8XT84HTYO4RkBGo9HF0ZTkgBHHt/WEuss/7yN9ntehaRNUe/hxTmXsB0
mOV2UXV7Iy9JFhDn0ztdVYAOzkhnHUe8oNLFPdMSi/akmJLdjn3689y9RiI4ZLqZWL2GBGyw/qOc
NGve1L0kHGkGQF0XW1/A3F0CnrKGwBqwj5c+ZPeOzgFb5fWbhSVzNjgvx1Esanjuhr7ydCd87lep
2jR98HxrYQmydB33l0F5WLivrT0nFE+j0bpwRg7YXTDkeRLtcC6/XVq/6wSEomF+QKKQTSaiSSZa
HKCAoZehxd6XTaZXAs345KzAlnZWDuhfTE4+4w+KDBlOPwzcWCH3xjIH3z/pXF/OMmdItkFmZoeW
znaKbn0Lyuv8XgVez7VcMN1O5lHimP6QmjtNMJtdV/aXbAeZncaI4hC3X+TKpVD5Sy43DShYM5hJ
2llpBfxSBcPiJzRoVeRZqs4qFuJ1VFD7lDt2xmCQyUb+gYDU9AaFaHk425WPlFlFltmiTZ+ghYcj
mCTw0m/+YZA9Yxn8C+LY1VJFmKQFHiqNK1WWPT8JnlBUXElQ9HgY8WRMMbaMgMV4GVh3s+0jkK7t
YngQqfqd2Wya8pEPqfTn997MgLIwoo+hGyQ5/HCkvHrSYFz330sen1A32SpMhdm+GSaMxSDd84nl
HqFnzib3UdO5s+CRfCQ2YNL1XLyu0VkHLutG3Y2hODjwkkDm9eP2AyRquWaiT8yQDW/FLNYbmXIM
y2i+mSjjSfG0FduBuiheJMMDYK39G7DumlBZU9vaT9JDqeMeS/OU5uG67Z0Z+rzBC6dx8yu2i+tv
lfmIt/SFaHUqEQTNblCIXCOxsLCmeDjhY8mU1VgjrwYYQYHv1J1wZEHtrVcg9Hr1ADb/MT753jsu
c51kFGGADSq5f8jy4FYiQNCd69eiMMa+wybEgYXNFvTQ7EBHrcN6L63Wiqp1exkvd3LA/MVFR6gA
+uCs+8IxxmD6GSeJCBY64NECjZPDKym2gBlQ6HBiCMhKVKI905XOLTjGLFiMpSk8RhQNCT/01+Dn
PEPLTKFpck58YqOlvnyqgkyjr+U3yq5A8uhGQunHAPiui/hKHQ094gOfVxo0bxBk++iwgORd21h0
i49zrYTcGqv24jGmRUBHaf3tG/vXWP0BJbQNHaBmfFQ4/Y/hZCF6ZQekwOcU6vFDbv4gFkM+vQKb
bxX8HBnxs7SwL3QpJUhKorPf/ba3TXJcNYSATEMikafg1sPduT66lCM0zob/4bSPd1Kw7AnR4Oon
qZRRSIGIWo2dtyaWb3PMCt4+gJIwCbJZoq6bL9k4dEJSx8GKz7DceetSssmsFsOeSEn4fhZJn3fu
WEW9JWp1aTGND4vy2/mgeh6kUeXe3oNaZSMOLzFlJ63wK6aRvI5d/Vw+4HxfuM8SwLp/lVUfE+Th
X9DC6/Lnz87GUyb+QkbE5XrjC37KLSV2pjdnMhEG8F8R7vh40NIxIPo6Q+p/Eb4i70STSdOIef5f
PQnsqP6Jq+pysGqrC8IfN3gVWlEolg9k2jNHq6evbQQHk7BUismT+WiprNDoRFEVnxHjjPbQ5jGz
5bTegFEL8i0CDSHO3bDvtHRmWDASer6xAvRcnST+vrS/Iohk1QhWLCIDSJSqdDsN6kI9eOE/2SXR
4Dt8q1U5fG6/Jzc9ZEuohn1oP9rlLbH/gxkmGTLnGF8ak5NRJB85TfKVEgad5qWALM9oRe5/VH55
mf+36FtaBdLtw1riwLOi9WUbZO2sMqSMPF4aPb6P2kLZWjzSd9UR2+f3IpCKLEwwyKMpkuPJmRvp
IE5YkZ2ZxKjA5ikTyXqr6aBKQdnTPkdtHDtdf32J7DiNwvUMRGnW+W/JVSMC1e5CuP2pR13Zrw+D
VeuBTAWYTNDelP/YvYsIFFsCKlPuMq9rr4Rxukg1KMdH3FIpGdH4fngCrURSfTfN1OEkmLwtZVtI
/qlgpMt4Hom9xJcisXH9xKFdTur3HIL9gckVyX1DKGo09VWJFqXwEAD5R2KsdcEWiPOJhReppF1x
DMMRbuG2AkhgxdqmJLY0OryjwvxBrsV6v8ihWu86OWzgGFgcRwm3Nc7x7Q5rz10TGQ6FkuHaQOlU
Etx1UTyq/yNv67W1L3rBDgtsNRgOZrQgq5ZtY9GcviAavcIIgr3c7+uVCrZT3mZCz9axibt54Scm
CBydF3Yuql1utjv0w3tjWH7mndQ4jT2ZPBnikjqGh5uC3IPa/wvvUM3VIKp3sRmbWjJ4hPgtGTby
loIgIUbjx+U13CnOehSDbpEqNAoADdPscQWCKCIXjN84sbkZP9PB4BPBxNy9VblZezOQCuC7Reuj
+zaCDY9Q/PSIffaeTiEymx6UmrmR7QuWXsqzydnXrmEbuEz0avdMRQ9uJzOii5CjHT2fQ52b4g81
/xuaX+EB7YNlyzkdhcfisMq4z8BvS4tCLrO0FDwS13SU1sXqr9CdCp2rPksE7/5nIiBKc7pCPWHe
S65Kd18n4NeCQHgFIUanHmyjlOYiVrLzpNGGe6Gd4XW/luyNP0BnqPxafbAdh5bpoUbWJPfVAHyY
eOmECvlVrHcqgRZFMKJciWGBPr0DL+2aWhwtnfX1KhcBZAjllg7v8y4yKg992I7lNn8ckqXdRWMZ
CzRdLPBIwVXXbwtY5ylpUCS/Q9MU8n8umP+ZvcFvKYCLee6eE5QC69pJBSlhGYc0R+CVd7hK2AA8
qAw6IpKw7X3+C1N/WXQBQs/QfiR6jOrSBwxdfwJFmu4KWD5dzSxRkktcHAMmjhVaE9j7v+fLWrLT
uV6DM2tyWeGwUlBGVRaRF7M+5tQQ4hPZnsZ+H2NRnMXlVuKOWtpWShgKjHsRXHePVLY8EDgL2yRu
UWoqrf3mcJfQxE0VNRt7pxHsQly4Hnpzf4Y+EjcXEG8bhhHZWvZMAAc075t0lx7eG1Id0VPcrc/z
YsEfOcHcJNAQj1bOqpjrwAka4R3Bo49PRb3eaCmq/8WQx+MNfO4fi6BlinLCQAFESeWbEh4ymBYe
9vdiqMW4GTh22WHmjUafFQsZfBCZUSgivBf/uWVg+jEbpBDb9/oZJnRMdloc/aSlF+gnPMlwHCaE
bb9LGzddw92/ywcow0KU55IBxmB4f5+AYLe2ANUTbb3xwMvDgPVPxcwq6az4zBvr7nknl3jIIxb5
vusbExMdfQiEcJ/sBgdJMvdlJlYz9xn8QUo11NCDRDyJKY4iUK4m+atLR6DZqL6M5xRhkDSuzTaI
SRt13fYfSYARVN6P5gcT3wMBmeJiKDeBkN9QdXRaHZpDgQLLCTWxmClaP04i7woRaAgoTy44vS8q
75T1rbgt+2hQlOwlGAdC5hEYHaytxv8OsroUeMwf277yc7CwFYIMMTdacqB1emYWRLxSEgzQgN4Z
5wFGB3QJQZTW+UU8x8b+vz7hTueEwViqIb7qEd3GfCCGa+ioRn/neE79ikgt5DMu0/uc2WfHXNXu
Plb1sPCW2pCUp7/ClWJUV7QXD3LSeBVuwffPt+CpmK9O9xTzzzqoaxs8Cyhs1Oxff1IZ8IE30nW7
huVgFglOkOQjfhBMmhADthVrL1NyXppUXcFAfPBBJqB60IWyYvfkxQaet/HXWDMbgqItqHLEYr2m
Qa8PF4SW6nWCWZl0L7jgDyvVTsm/9P2c14c18YzinYkF1WNFQhJbuCMJNUVpihH7DV9rBhHY4KKK
/V2HTpSR7H4d36rBDNoag1o12f+4YpnKQYURFDR2MQi+OsNjLgzl89u28EgQ/vUb1nXUO+pJffu5
cmwpoh9mcYl2z28cyPthfN5N8GeubIq0GZ3oiw8gvdKFOAZkdphlRuXQdv0HXnmE00JRX4T6gEAV
P5QWBLu/HWcBeU3UDxhMqU1Bl7Fvq03hn/AjK13agX+rLhWBMXxejPD1+YCaipJwGKq4Zg1poOa/
KJDoze0VX91UNm+GxJem9f/BQEPAOSTi8DlmSsiHBjHA+o7jw05sNfoJZyhgC4RCwLMGZaCMRwiS
f7s43V1aAnuPAIfcC4Vo9thfISpm4a3BZoRGyWboIJuIoNdCn2FmMHG/uJoVbfN58faLyMkFJ7f2
RiPWSRg7vA0ba0ZiY4G3A7p1+/D1b7vpQZOAvR/UdplsTuLwP/aXh0IN/g53bQS2GuLOPtgX+ZiG
1I4wyzE3nuSOlG3OIpLqawAjSCOs8SrzaeqyvB7EI+tYrPw8pcmZ+zfv0gL2c8I1xr/Y1JC8jo/q
SyDYP78irJTbC3xjNECeSB8Ej6SrBKyrtww3o3LtRRprHnDHo07iBsX8pO2l0DoC7E5DQNFggE2d
FvSg9SDPcqovOcfi3IG9VD+ep9QFO6ZiZ66DmTCl109WcSiADMg7GvMbVVm0vLfcLePf2X8C8bWR
83rC1zlForxZtWdGhbNFPDJpJejn2juyb7ZBNSr1mbdF0lAvlzlHNFgEjAq3VWxIR6d5tP2VaL2w
KiPvj4Q0UIpmf2GNCxUC2WwWPvy2M2gINSd1fyDUn52aJGj7EKpe5io8AhejrQ+TbCArprhzWpkP
ZfzXhQiJqaiwQKPootw9Ut6lEGHrO5pxbnAgx4ZuxJxsBf0vuLeGAQoMX9DDOwfhHsEv6RxTjtIl
8dVMUJbW3mCcYMyGnF9z/vo/MknFPogJq7xwJ4v6ORBfjYzA4YS0UjS0LQi6uHRu/V8D5TwgURa0
mkMt0a2DjIYoPl+V+xsu00f3i+eATmgomrzvmgp+f5HaKhbIrLTE07ke30/g2arljnRA3Vs6vj+O
V9VEcJTllZsSqAN79MAg2qKpHTT54ZkIw2PShE939CSOx9Km3O2wyCs/GHpS3bemLb4LLJw8lxWQ
cdOyrGTzzzNJrgpEnrAuUaRo3gJp1QQVCUoEnI25V3rXKsiIqmkBXu0NFWyGz/pRf2/3KtzAf/TP
I0jE7ysVpew0RXnmrhSYOnzQYVH9kSGJFjE1IrTZ70zYPd4oA+tTzys/6OQqDPn6i27a5ucqmZGK
M31g6wZm1RGpWLZ5u0LPmozPWH9O1Fm0Jz3zv3iBxLl044lfNzHSwn3VPhMwpaQi2+7V5h06A1rX
VYj9V4Zm0xblx1S4hd9s8aB7HtixFzYCioZRIONSnpcL4pTwg+VELtKQfK4jU5zs233QExtuaKhN
wofBCR8wUVx7M+BUaepOBdDDW9Vg+D2Euu5ht91kntOYM3HkbkAUC1bvbnXt5ePa/XTWtRDAUDxD
zc++wd20JHmNDgD5mPflqUxTMi8sGYfWUTMcPiUhOsfjtNr1qOEaz1FWULg2C4CFM7M10h4k+ITR
f3fEvx8E98ScHCaD+Ad6xPgoDdPlOrYJ1v8nW/sq1cbuH3tYcVB+R7Xlxtln1UlyZPkmJMK4+c5n
n3ovd7tkyucvsddm8QWA+8se/9AChzLIM8a+sX8RyHycWvOaraoXAUAlOWsdqmLvaIxlOfeD9JO1
A8Rn5wupdEhVQpcqiSOhjDEtVH0oVF0t5UBSWWb9RhxxdUwxE+AmatZdd44KQ5GjqQaVLhTQJZwO
eY4jQkKBEUz/Ynubi7vqF0sGYJedk2+dhSTbbRbbhwNJj8vcDh6h5yJS3VD2hJft7iBWO6OVZmcG
hlMZO6cM4pQT/l2PieMmx5ZyjDo3nncjyXBavj8QPaeGwVTQOIhVZ7uXh0vp3kqRuMkVBbU7q7y0
9fpiZ0wN+A96wKjPsrNtv4/mczN9Skw0J7ZBXkdfXAw/qGQFsf0OpZlVppsFh1vUgVCgrYDSMQqM
2RmhWOZPJxpW6fA6Q4YwJIfnesJmZWqW0bgm2MOf4vx21cVn5LOdZr8/Mr7Q9vFkahpe1eEpmdIy
Pr4MsFK/VMUD7V8gWSlzatSNPYUthKA0vqS/7GhBG1RrdsDVu0Yko1lrn49ujvhg7JFC4zXTDyw+
qm5AQlmMsNgzQMckpm1tTcnD7FdSrGJj9oLO+VZWD6DM0v6/qWmnO1j2omt/NPQG9iJG29S2jcxb
fb5JG4xvDrfybYnUTd/8UiAMzEA01HwEUa74G2tUZKtxRQ0hdVp1aKT9B4iPKT0S5B78dHIX1xpy
pfFWJjoSu71OO/1wPBbOHAXu2KhjCcTUXTGKZkS9a3fzYVVwffIGp+gR89cId3Q3YoOxJyXbY4UP
Is3n/wpssecCqwpvLAzaE0kUZahFjCZxtOlsEqUPGeTw5mIIlvtb3ZCqaMnzBfHN6Hkd43/mRCFx
+gzcwRoFV1Q9q0zyHyd81LJW6LrhkRPoCJ4cEQoa3/GcBVsFRlNNuKQXBEP621xbO/DmN4RQ+sX7
JQ9moezXdRUcIbemsCvCAeM9IU/qr+pEJqNzamRlpEunc1wqMYFD8zjB5/viR1vYagU2jL/1BZdi
DPEqPZFR79FyyW28C+eYFZj4l5m0YfUoIr9zs8r2lbm7PJrt26zBOM9sFcVIpvrG8TxVwoSY29Za
aHc7Y+Nitn9KOgvZkhs9Tc7VbGp01GtItio1OzJFzzypKY5Y8qWxRLdcxpzwSJzTTFi6VxSnwxky
wB3SHn5xaKA5foMwXPPrdC5JpAzrSoqIpRzi3dCxQgVp584Fnm7p6Q2snoU8e0Gm0HRYqYTnZLV3
RnOzLPFM72dH0S0AWjXQNS5NGkSvL7M4SmhySQlB5OZyZfXneCLpn8+PNj4Bn1XMDvqgqMM97ifS
L3VjtmdDq1jH8RQN1waT4AvfFNUJR4a2IjUN7tv7AkmUfqST16ohYU6EKQP7vtBKnVJgW/WesEl6
erQEyqbSmjd64r6hNXliv/UJov0w1t8BNXfn6e6WBABhg2j5pj7ghBV+b4/yT1C+zxq5vfmiza+0
WOYE4fvjoU75fgqKva1ELTG5pfmwfFEkNPB96xd12FZVu+wbKY6u2CavuricnUma5t4/2WSVyayp
UjZRXXMmSicELCdvuoGNQRLjZI5VipHmp26izuIN1qVq5oPhfmkxrgehd/HoBrDGEG3pzfFkJhAY
IyGJupdEb3JNKucAVX8IVu0u3vRsBfpoNiceR9obl5eL2/++aTrEwaINwJhUjEbp9vYp+MTeEprr
1iCn6hVqObOfVIKPtCEhsZj+xHLcYaKvtsTDDztZfpVwBL83Py5dx48uAzb+FWT9VBUZk/Zm/G6I
/FN58WZmKl/pcBHLuezKh5BoRs8qKmEnkko1exjg7DhS124z/pPJLLUewhsCndMK15kOH54u5f8p
EnpflM+o2u2z4usJDL3DmP6AVXDG+QPjr8oIQyXkHUGbtusiPIfNKozCnHN0mofd6aosF2hg6C0K
VPQemTGn1zRI1syxJMgix9IO7jc31mxU7BK81BykGPdeyuf9II3uplmvbzrTcfC9Qc/q7LpeFtdn
VFGedJP4Xr2LKXs6sbcmYyn/h8lh72SeFoLFEjRi39/mjIHVrseWuSWuJ6iX9E+XWBNMBntLpdB/
bJFwOuweNMd9rE1shr6wEMj0nIctu+usFk/fnpF02sRbP5rblgIyUrhHd6otIAKWbPHoiULTgFpN
NJOlKsZ8h3v+MvZ31Cu6Takar/N2fbeWMQntYyzlsZOywoLbo9K052guK1g10jJj1urBo+PLmEuj
7xetBSjDb46oCQ1glKA4srv2pVAqwQHGtkfxnJAG2IF9kRQXc3mQGJB1r2q3vUWf1zLdEg2072d4
aMzZ6opET5Gg4X6p+7iNRJbdhKs/1JPRq1Jf1wmn+MhNAT2f2hDl+XEEKo1cfwRI2Oc0Gn7/hM/w
Pe9RwljfugL769wcTbygjzUcQ9zUqc6IkYTZVYmD0v1bbiYWQE285iZBetLPctGWm4IM4lQ0Oz+V
2tFCvSt6ILPqypVMz/di5XcA7JjQWGwwspxNWbY10TrjCBTbcum421umBPCKbMP68E5IRdbi5FId
cK7jCHoCGlhg65zWonktXGJo76di5xCXEkvNY9oxhesmyrLt55uhiVl/+olHzfEGV7qqI7KoaRdO
l9VZCkv4wuQrKGaBxQriux+B8WpwYOmdF8/xApU7HfwVemFTOUbw4oos5ZXwcnzUEQj4uPmJHBB5
g1Jwk61V55hjQDJ/kxZ29mp/0GV9yCRFoe5CHdWzqWKkogCfBKmQy+Sue2bRXaaSzZBzU2AN6uAl
gXhz6REBi4j9GQljq42uv/R2SgVYBRxgi7y0be21D8UqWp+iK/pJjAZ8tbBsSipLT9FiC5/sM4xL
nYGwffbTyYKI5Bxcjq8Etz5fkXw57HgrI58E/om8XxUJsnL4q0SmLN7mPsdXcbjB29ZD9+Ghfi5i
F+TMuoCe+80C202VnzXseUolroAj3ThqX0avQkWVDbiQ7HIaJWJMK7RrpB9v0XXASruLLgTJ22by
N9zgr7Ro468wi7zWNan6jBgYV8PjiXJLNpcyBm8VjQeSjINvqleRv/lcS+Kj92TChu2NV06x6HVE
ucyGSpMgycMbZrtlBSA9LdFR4zoo/xD8vijkuMh5Dckw8OhG1BCiU3W5irYR9j3rEcv+BSw574K1
oLbSOCjwYV115roTQrzASIG4qQcKb3O9KvX5pgXGDRpE/VS0FxEbk6hQBZC8omF9lq25itYGvtor
Y5FHUMIVLh+M48mjhxCQQt9rIurZvgIgWXH9bA2kuun6qxi+uZdqJfDCbyXdgqDUV4bT9v3Y4ZEm
otVvBAit86WcucuPqEKji3F9PdV9rUjpgrfUJWusPGKHAHZapW8Ttxd8kbX3SB3d+VmFvRThpkjd
OcYy9F+a5iOcxruyrDO7oi7Z6YPHvssmXdmyOYwOc389UAX6IocDR+p0bH8NpSZMx1Mlh88xv7YO
z53Wd45UEd4M6AvEybuvGCSB1ROjhWlZcpgEG4K7idIn+itN6Mg/8JOXcL9jiZjl/ZW80IaFmWjG
jcyURr7uCLjkJSspYjo45qJPo//7gY0NV1OkZF+WSB2s2bIufy8gRfHtyq5/sHOQnS5ZFpIEl0/0
pRHWpfCty5sBJVsiWaLXssLIWvzjN3I86kXIIxmaGKus0vOQOOOELrgAsk0P+nSBYh01H7H8rzkM
C7RJCZbMNSk3n14t7VwsIF6zzJ7XYRAM2OTR0/QmHEmbVgHfQM6hK2S/PgPyhaKp70zWqbvXvidm
dwmCmHN7j0a/lhCuCZ+xqOxTsgziZmbPqZEBHalx2JOPKba56CxJRoDE1AvcIgx18T9mHjDfF3zx
vrsBBFmtGI2eJA0tgMQXDO/GwKqolxPJBamt7KsNce16UcpFphyJiYaxN5cez+7MEoXhdY9J1VNt
WfegFOiqLYUQ6fUxAKdjfjLnvssl9COtHxkJX0RzGThQwN84wvC1D3Brvx52L1YrTF/Mofeko4li
5SBz6ftZRA6h0yTNs3xfZifDxqchiffqlRYu6ybTyuN0htVTu8kHUPxey06fX5XuAr9zuujBHABH
TbhEIJkWe0gpKg9aOKH1Yaq1dVT98fVDg7fSqXxf0h3jLnQnIDhsHDnJJl7fiqKYS21WjsvpJAEU
AVDA1RaQWKqJW0lGORPoPfGBYFUC8gFDXrGChM3ZqMWR670iswWwL6oREul44LB8y7sf/Wr4mFkK
6nG+/bFm/SYh5jWdOAtNZDSDlYB84Badq5YwaivulxOnVJPYbq3iMnB4VAzXXnG0lLyopEivdn1E
cfm0AWeGKEVO/a5rhkUBgdBj8GgLyV5pye9534P/BRVa2XGJoJWauMnreQPWrn2b49qK9PC/iZQM
ch5nIWhIKMjc2eu568OUhodYGe0TF4WVfzFjgGY8J0y4HEqxporJm9VZSRGqvOlBwkYEoKBHvFRm
+KE73dNDtcCHUyxfMjdyU08c64Jn8gF7N7mLqW6/2oZqPf8PLlGKi8VT2lusuvU8Q0z+Rz+RPksl
zaIleOasbOLhYe/7DQA+rMYcjWQYR9e+W2nQjdRlpz4pg6jZY1T3LdjewRoi12J5/t0zCqSr063K
L08Lxv5EHIt+LlzrTQ0wu7mB3+rW+ysNC81lDo5IBsvwObrYlqtEghQoX71sQZqVJYdqOaICbpns
uzeWkEsLQzW0jo8MjVhnR7k3Ltpe054afh4RogRRGSdXJEDdGtGHLwNZ1qUByAHIc+3EYI8TeReV
/PJ3RBsAc55H7Jh3m5RY+rKMiCID8qCVXkcx8ZD67teRMP4QwV34cYRd9FPZpjafm1KPjEgR8Eb7
Hml7b6P4B9rxHjd0JyzQr7Qm5CGVl0BW3F0QsF7YYXfK6tkA56/wN1CB63Mv9sirKwq8CHOs5XXl
2f6LYtMrjax+Gj7ecoO+ppzzNpXlZgBzQxai2NsarfE+qqt8KXD2JRmzNmnJMLh/1aJMhIKZH9LO
PEBhU5RGR0jxa5LOQMMQuza3DXOqGX6k5J5U6o6PE+1geEZCaTm6IQzd4zGOM8+FlhKXemmFnQ8f
mOqjJt4IIPAg/Bcpw/W7TfzKqPo08Ka5dYLOcE93dpP7VpjQuVZll1byuYEqLFh+jFQXLtTtRPbg
SYOttFr6PfxyFC8eMQEGQsnKD1eMoe2DWfZavRbFcJL6cbOgGb1gnXxaTzYTSZPOnaIPFDwZ0F11
UuO20/iv+zslemugFhDVZl8XuqyUtE4Zgd1lpTMUsbG5IdFzbpiHIOo/juNeX0cE9ttbpkER6Q9X
UF1P3N5Mk+fVEjDtMk5GhITIG0oG8HBevgM56Ud/rvy+9pXFk+mqhmp1hQUMSM2XxPxvHMr5qo+d
m/agGZEEAV+2WG/lK2pXy6ND8YdSi2ocbYoJ35RuvYuCvFmN6YcjZfjerAm8q6pE30FsubNejVfn
fBdkK/rJYWJFieG/dxw1pauuHtOMNuNUJxGxlFmOjVYVdsoTG9lG1B+0XYN94LibB3OwoyFYEGWr
pOQqtSBRwsMEFIHf84jCNQzeE6AVQEA9W4fp2f3JcRdOsbypEAhskq06rbR+iFD9hcdu5ImehOP8
VFs59DiNpK6xy67lgyaNUt+tCSmz57rcQNaoebpdcQ1bUrLi7LizlqqUq9+uSzsq8EKB4CIb9a81
B2M3hA8ii2XF4kHzo4yQj177vqfStdOBrFWseTO6iJoS3m+6kTH8D6gDegtURbcRRPLuJl6BxMOY
TPnyZKojM6mOanZSWk4ZPg1NlJ4Oop8x0Pocb1s+JNXh0nD0U5aNVXbGcuvOhp6bUEdL6x6eP17M
2NhWqJ7yzqkSsp6lUTMPDv+LMcN2W6ISTg/u+ahmCHKOC/IP2pK559LFWlIRB+G48cdD0iezV5om
5ZGUHQtQ2va/D6QKTEScYEEBGCwZekEGeZ3j8qw4yAu/nmZJmvS5K3dIoEULXvw3X13uPZqud/uS
Zl9xBnOXo+5CQmXBvCqORz1oaBbIM8zLXlnUGAiFBVLndP/ADA3y9rmIpj5/j5CuOBeKfa0YibNq
svK+tBoLw6fuRGRHlpai39CMO8wGVhse6r47qgxzcanc5gbVnygfCDLs49COqfmUg1SBcOJiBYEh
zBHEfw0c1IbpPUXSsQLJ79cQw7rM5HCc3nBAgO7Hct+Fv3eYcsxQNA5ILxtGwfBX+GoStpnAgaNu
6QYU32heXNop4l+dM1DI9FpxircdpIcjv1diLqOdohokzMadVk/LrKvaCprMfSm4exoyeMjjYFDO
DM4YViUPL94+yumLTLl2MiaRl3QEylhJ7T4Hvvp4CKWVeawkqNK04Yhe2006ZJV+Usakdx/HAFPk
cDgyl057Jg2Q+Z6aOLUJrDYkGraGK56NRVOHl1l+1d0f6OLrFN0D/gwFTdDCCo1Brxxt2rDt3uor
KXZoQKS2V1Y+xk9fBURsM9sJoSiUPzTeCO/xJXMg3dO5zvLK+Vulh/R684CTpYScDNoQsCMvL6RZ
Z19i/PW4z7jt/hwl6egUa5rsyoPZJImzces40yEAo2iqpxYKc5r47EfZrWZs+/n+oOgTyORvpycy
xvWeOYS1+hhHDWpkk25g1AB6Kb7qMJXG1O1A3Uss4tb5EwCzOD9TiWxbmAsdCeNgdMbP+M6N9OWS
DBXroc1MMXV7maxtRObJf8QmFdNRN3B7FpSJk34M0VXgMiHz46pw6mGY0htVTWTtmC3GDrQQrlvT
h2xvOBL3/padsLpEHQJgyxpUObqnOhGj6va9LwHyrQ615YVVQEYIVW9de29PqxNrgA3uI9d0k9Nk
IuSe71vKFLAWQ272ILk9v4JsuQn4spYeSfRhJQNThjUezhgDiKNLbDc5vsnz/Kdpa+H56G/bgc0B
P8MWixNX8+cv9wypESgj2seyRt7+SFIwTLrrAAd736+tKtFCbYEWTh5hzyVbghJ1C/G6Js6st5Si
k9MX8vK3EvqDYFJqIKb5+N5YoLFKWxiKfSMwL+btzBg7TfS7jfxgTQXKh5sWB9ZrLnHB9bmnwq3B
dVc6eig4h1juJa4YzCS9DBbzn8A9WAu+ZEk0kUaUXI5R43iLIR1OAzuUf/645P/8bOdrjffP36kR
eifRWV14BE1Qc3Co0mmjgbGV9J0D+0YHeiv/EuYtiJXNuIb2B5NaViRYsMRTlJPUrih9MTxjiLGx
vBX6F8mqGvjUnb6jpud+qTR0sWas6o/eF8JWMHnOlU4gJiYiAHro6drrTdxreXGLpozrLnby8Opv
2cm73u2qQI+AWGxTgigFq/w6/RwbbyEQT4Unx9GFhrXisiM2x3G9v8PnsgVVbcvk2AeqKhdZ4Z2k
qmaYDKY1NyAyTrIlpmuJNSkNJ3VhoNmWS484We86bELX4BdTJsGztYepDUfzYi82miHCPjbWiYkW
URW1DFUehrWBs900xM8gL3naLVIFEWUBwlsdrMShUmEIkJ3kGg5yWsDVJIuL885ZMNWgB4qlw55s
kdmUyOKtcTJZs8ypCTA2it4BwrXKJQbUYQ2PTT7yWdvumFxPESwTrHuz9Q2bdx57SNqxOMtaAH3H
gc+uThdGQSNBGRYH/lsO7mrAE5Lhk0q9oQzxKBpXShQc38MVKGDKaxUQuOvJQk9qUwYfpHe0JKM/
KGSjdpL+6gFSJ2QBNwjeCS3UxglAzwE9j7BBv/O6NXqBWtrHkrW1wtmmOiGYJTgVdyzqaGC3jKsx
y6nqieWcAa0mzZnsI1AxDRM+qzTnfIswD0lFtreg4cIgTB1L/wZp+nwxgmLKnqmtRPsHq18Ek9ho
b7JqO+cK/92YDeW8Zlmw9UiraQGjpZJNvQfGzatd4GwmMI1E8hZ8xDBEvnQMEdieXVWkeZBOXueS
kaPzyxV5v+Z91ZFwJlw3pNVjkUhFVqJIg8HAftrWdH7WpNrxi/pcKMeIMEkC9LzuxN9W8OYay569
d7OIZU5eXfOBtWAnmzMGEQS4+Bi/7BFEgnypE3tggrAgliqlVPFc0OIjvb6tL8+WUyLlh0/Jfo2Q
E+Yj1/0tHykG5/w5MR+S6qCYLKNdYi9kmqgEphLSwmZz4kvDvMgYRW7WQ40JYBI/1Io1Wsk4B+vF
TldIfoDqWXtCsrx0VIp3hfE3jYGKcIWyFJHF1UrSTTwuzAZetGE5RbPjdkYiNMCC7oPqIKuwdGKz
IyNjdWOFyHXbHUAW4JnvncHP0fZVWcGG657oMaRGpBOghpstEnM/jkqld7lPjlRcj8hlv1hS38nz
P2w0p+QqOi3Crp/Ym/F1IbkSQ5DVe2n7gTbIE/1WUlDH4KfevzL6Y2+1x3VazKQk+jPJhIq0oueg
Fr7c4RP1L7XxepLbKBMO5DxJB5wV0fkI3kBU5oBY1JwzNRJGnN3K1nad+K0+XxH8ns09r26HYuSF
k21TNg1iGeL329mhpvh7XJhqZgrqAGeR+04DN3wTDIN+1tQHDtMRPhvlMyeRse97zeCrL73CemFo
E7GNePk9E7puYUMneUBzS7FBp7FxkfruWNuxLJI34+MA8K5hgc0/u8MCMOZfKbQIffK2gS+r7P2p
s/WPYS6XAMnYk67e9WPl055hhiSLpL3VvIbd4sRzHcKaHJMuRdv3N8NCM8MicG7njWOnmbOOpwIE
x2GAXwzvduZU/5ug/qomt1iAJMa319BfopG24Gatv7AQ1rkLXCgweFbrOeHccorUYWj65+1rBDGp
VyeZ1iYNHopCk/b1AtW2FJoP1tuRZ0LUkqwN7DAfp+Jd1dhCY9ziJjQYExArNqczwaw5fs4IjRMg
06OZNc5PRc5F7hyyN0SluQEaFissdjbWPcXnkfEkLsXfeovhaRnxAXsOBAFWcOi29aVFfdo3VTgq
1rFUVBeoC6kdMYwAUZKDgLU1c/WAkzCOY9z9uJUNfBlgb1E3RCPLVU+YNjhSnaNAvkwDlBr4XmRo
8AyzpytAWbufErmXxdfxAsyJl1ErEFr5LxjllAiF0HDa/wjJoihJ5IiUfg0HnJJDtR0ydJ8ngDRI
c+X+KonvdZ051Jr46ZigfYED6U26L6RHUlC0jqhm7N7ReLd0bZHESfU+tcAdUt6uk9akfZbOGnfC
Yw9MuTjFei2pZkzWDzexg1P/z6tRDq7tZ6HXlr4yDe9qJLmQh4pBTLJykg8XXjIvL1kTSRY758hJ
rMb3KmnlSShmpsHussroatdCcd6AkMltEkq0HBN1al1Wh9fnufsi6MWWK7Hfaa1WXI5AkNKE/qZt
Vamo/mBmdhfLp07po7OCv7KGe/Dwa9kqd68lVsuo3oMCeWQ4ApkcyR3mvVaZAmo+MaqF1mcxuE2k
vHMividLGToXqtzqLbNKFB7bsK1R/DwU1CYrCkW7STnO3RbYbQjex6+kAU+BS9TIiGOPFfVhhMtF
JTnqmbjgCeQ/5pB/FpME3zp39gD3L2eAX3uRfo7gSUD/djHpYpVBbyKEzkRISZms4eA/Luwy+7Cd
yKISqy3CVaGU9df1/Zb5a8cm6wxVsmSfnVCkUagejPpVGUq8+yBT5VABGPT8rQdejDFkBNcyb6hG
pHKu4rmglcHH1PlJdPGuOF8objk3p3onHYJJ9XcIqbijn3Gl4t8rW/dlnWRNk9sqWGUa4To+oefe
c7puirDKEO8Pp/N/QexPPYqpmLRRW6KY/mXTrATCmWvxy0AAHTWurEzI8DlMRJ+Mrn/BVLuePRCv
QLTLNggx0Qnott/3HDkthwmr7UGAdeMOrzCOvx7Ka8RB0UDn7raS+QHasaHj8T2JOEo+aFTAikfV
YFp//+46c4dSkdADhnh5bmkabZ39RYuYc/jvdLFjbw+pCOd0j2/NMCHVdOXCiGDPs9OnFpKYBsC8
y/C54WjWXpkedujOFmqv1KsIDLXZZogafyAv+mei2XUCNaDnlSZbsPvv4H1fzrIuXMnigtM2CIjf
mRk19XamK+qwhV2i/RJa3h6uhNp7vsxK3DMRbLNoY5L9mooPiU9UduK7PIvAhLTCDcYM3q0UE9vW
PchFOXOdzCo834FY9N8Z3t7EZHo5aI65eSlzCSCFTzb86XKWEBJqhvupgyRjqDLE7ZvC9OydzEIr
ITU+DKk+CIfhsl9D5smev/bSMDdMCrfmarpS6IwgzqXW8hV1ddY9qD1XVolkSMN40necN3Qrmfd2
FKDf9knHYXytZ9Y2D2bv+VUw8ZehAwbRT/5Y1NZkgY0fVSd1tIOijUERPdUSYtmhAOfW8xAYXYEV
O2vnv6CQjzQbBR+scGM30eZNni6SpFCOC+wXFEkxx8/Ycu5B0PrPTT3XF3c+DQ43sicfjUhVJsLR
rL9xjZbdTelh5FV5GK8PhjIziz3QiS2TNwHqzgB+uPIOi0xAEJj+Rye8u87YM4NQHlkmAb3t+umb
xeX5I8rfQOr8YpAwjjjz9ZO31kKuftk6mPhy5PaeRx1TXKA1qfqfTKQZ7Vzr4dh5QWPwComloSfz
NzqE6Zth3YZ5hS0dyFkGXadWurA4IJxP/oyZBdurqDe9Zn3DrRd5N9b0clx8vy0ZAAOVD+xJFKf6
5/ufXFjMABmdZIlYp0dbbXVGNOXwQxBrdYkFA2blx+QDQZra0l6v4pvdckEjRzB1bydDQID4yMn4
NeCpzastTBjGoqbvNUIHs8GaugtHIQ+HnuubH9xp3YJrwTBJtSei73qPKWVlq/WlE4OxZR5glS8u
jd7QtVQlazPj6Tm6CkuKn37vCyOP+Omot5LKGYP874CvPqUoV5lE3OyI/ksarWab8H7xOYtN8Mqz
BnzN31gjafLjdUbFsJw8ILThxJtgwaSezCofA3H8qr0qkCH2R3w0Pe/36QM5znoLksIKDqDo0LTX
szhsrKpZI+gbSqM6L78MyvQYPIOCO/c8ZOYdUciORKDfOyrjs/5MPrFeOc7BF0P6hfZzJo3awmpD
qx+iLMbPZ1VF0s7CP7EBj4wfE8OwKdabLZpbSBNVWUE5Q91kdB2mlbY1spWXY0hxuIhpPTxYx5qq
CRGANK4tdFBCfgb0fk+A+QeHOQ9xUSGdrgzOLWId6WS++MaTTVUBTo/rjXYh+1yKQKhxS276dhMm
MufFKWFhETasU7F/h4AeaBtYA1Plgy3HqEHHrFBrG41AKfiGEo5AKhfuqMEO6q9jR8Q75i0R2PPZ
RIPmqgTn5yF8tbtTU1CPeX3IoU3CSwMxo+CdCAx1EzsbddNt8rqcfpgDvAPRurO+tz16Pm4e/Fjt
ChauAQsDcGwB/ZaEmMjdtG+CfjXrPxRaZR9HvU1UvtVHlK16zIfD2RXw4Zn0wlHIfa+vY/SyyC4z
vPVgYqrlITASH3DUOQw7YetEaDFuwy/jprYQUp9rIGHccMz+MeF3F4RqCDgAIityt5DFJztdX/sz
VL8Kks8KmBWYlDocpW2N0VbC2MoaANKnXL2x3276+iIuh+cacijFJH4jR79kHUmts4a6tWrxE0Ye
0Cti7XG04PStZQR1NmMZmBztwJEv3GtFfCQAU7aNac3fcv0jcrFZmPgidELsBCKvFyPiACZCCeuq
zTPu40UN0Os7rXuPs7Gr6lhgKLILr/kuOxIGJtGClbgJW3q/VuAjT45/4ZyrUcAR+VyBPqH6SIBK
Lzji0hAczP0/Uymnuo0TlF9ojikY/YsLYNDgaKCsDOm4zUbSI9yVcJCAq7CfAqAJf0ZAyzN792x6
Pqg8OukEnvzjktq9lB5b98Ku+J2xQBUF52jyDarkb/7etvh/WrXmyfXRKJkxqi19uvpUmUu77NKD
8vdG4Plm+6LcWPhSM+bZ3eFt2XkDnc8g6jP8B5UvreRPy7jj43BQo5Bdbv+VfKWcirwJuHF5oREd
NXZX2b2xmLOkADXnErNPxzqo2AHk6rxVa5zCbLn0I7IswUOVCFIMxSJDl5UyN1iey8g72aCvOPmn
6aQGqYcpZD8ZgfihpTSc/nozp8ZlEIpJPp7QBtUA2Xgpa4lNZt+nrAm2rxrtpoA7HeTGEW3FXs5c
Xc6GZIST4zPfsYgdC51LrrDc8xHWCA3kU1aDwFB52DbepAwjta6Nzqo0HIVu+BYmzAPJdS+l/uKS
GPgG+yBcVhttJ2OuteFDn+5+PQcYewiglGJtgeLxWLYlzwzsGp3XctXkluaYCuAdaU+zh20FAJST
SNPkB4z1MVVF829djGdO3iKlufv2CU7oAdsO3Q/2wIPYvBXBxNapobefjJ/xb+2ElPiTc+2g9/0L
NtxMqUnXkOXbZDySancxKCDum2d8XDjNNCHCvT8Z8HDQ82gwD5RMtrYjEsBdV/9dTFDYeyQcHgnk
HckbCbXGaOzWRoWkXEmDizq+BASe7r33/kQQ9GcjXduxqxQjP6nl5mJ1D15pmbE6YFEBQELWD0cd
xRK/6RSEMuAq4hy5ojXGe/07V18vSVnph7mGiFfJN4Esu8GH9HW+P9cwBxxkWrsBPXFr92rH5g+H
BgbzQES2yi3rZvJlTWvIUyP7OwuCFJrRcG8pvR1vdEcxXke8La6lBLKnadwTaMeqocBKQCeuugCE
e10Gv/2fAfGG8gF3jr6SOi2XzHukpb6ypyQO8lNomuloSiuq/FrxcozGzt+2aYuvcS/BhmdEFXYF
P1SdZPZgsOPbYkWfF0jhCIXZOYqoI7wDqrM4NgtbaxAL2SAqKMbipWLAHfApdPUqUljUG+lehjHw
hzpV+vPoCSO3HbX4NtmgkK0MLZgGLs1u7IgMDGdU1wRNSrQcXH0/TUQZUOTfRQ5QU/K4wdIhoHeS
hIWfHdFtS7zkd8W31jHjozbbSiOFndm7NyUicbAIpeJoncpVnymx7ljVkldI6sApwOw6QWFkEt5j
9TUvo9pId8isHVpsMYBNPTWTscgswp+zDAGz9F7mWveQfEBuRvq25fA4jI/g7UHLFFsLRLxaxIgk
NA2/Za0THNLkLcgIqC22QhKHblP3XlSFJudU0/VtMElfND5/FCkd65Ec3sek812d02OUaD8kyjdo
pzdHWugk5b8h7MvhAZYUChj5CpcHLfp+nxf3MBzPp7bWjhRvs9Rv/7dg1yXi92W6XSWHTofvUOvI
9OuJ96bAoTklE5LUJtfkCEGuvzw4FOms+28YPa2XhcugBGfidxDYB4CzxtQ5U6mHjLgn8du6ebkx
tR9lgRtWGkw4Hi0Mhl02MSoHMs45rlVcIQYcOkWa0ycA+2dDktwESWJQrv3aHZNvirMXSwS5waAc
AOPG46tPTo67cEJHUVcWnwaRTFAUpfARdsG/rv8UYEqNiSX+yjm90VlJjlfDJAZ6u2vyik8EbALw
X9deVZJvG0mYrSPXJ0DQiNOWYPIanaEBje/ts5GpKSWYf2JTR9ZiJ5fwIUsQ1umiFztQ8eeEelYy
9Ho/SMXLb7TRv5BF1Hu6ZaQZcthG/EPL/gkhfw5WTRG+nhLBHOWjkJZiZQVnE5ihgQtCBf6xHobI
3/iPAGkRzZPZfeVMEXlEkCa3MS0YVa4Z3mhqSfgyTsjzFMmVG08+LBHY4FcdRchrOAE+SCZOgdlQ
x/nLY/8sBegiWB9A/HfXltZsx69Cg7Evtrc9gN1N5FHYCdxPKrvGLUKdcdwxuBQMzBC1AJ3XIkFE
qFe6qPNYoltQnq7Brme4L16GDWW06l+Y1UfiHbZ2LPEAaoVFor4uNQ4TaAUnVq3rJsA/OIzFiDKP
lBAR5eBGRDf3Q2IkhcbNBUJR6ecY2eh3jk1zfFuVPs9olY21jlJsMPVWrlABHABJfGTJGOjW0v3m
JyFa0hpJTlxzElCrCbuDMYZZgCY8K7dBd67+08cnzkIROUD9jyC26K5AEVnIupQBDaAYX1UuFoWA
yRVOloDpRRxNT1eZSybn4avWkHR7LpR8ynHgrY6ow9NYqbuWJ9RPZTuYy6HEqOxYRkxCEvXTsb7z
qTbbnveKxafofJ6AjaQUXXwbzKQkkdQWIMFDkvm85cgZdUF6hX/o113tojbYTkfpdTVLr8wAfIoz
QPC0gwm48LBHNAPiKWAvahQazU7mzhoBB7yVbQyIKwuq5SliSs/GPKNXWiP/h7tnSAqeu6tKIZFe
A20Yp0jZxbgqWEfggrYOVKER0r3m69kxdmz+6HDBN84qtlsNTUhd7crD6o4JiWTgpo25Wz+/pcjD
NcgaYMTaS+HlA0sqC4Fz6+lVc3x4l5FI9MC3DvOYsvrMjnsB1tjgU73QrB/S0YZEhqEONTpheXAA
mSk3xfD8mX8nUzXNnhU4tETNE7vWoJtDCqPsv4PUy/svJ2pJVZwgcvWQxiDeTB8cTwf7G4LwG5a5
UVV1ueszPGkBY8hbq6tn8+rFNF1V2RM//y1k4xE1e4nlpgY7Zz3zrbew9EZbNcwOzVzDHmh9rx2M
RPdRqujTCOcCUX6iFR9PltjGxtsGP3W7Qsl09VfGpdtsVHJceZMEOxvuULYj6XMtF165ff4avo34
OZN5dN0CAXqeajCsqWfHiT7icUssCyRMZLPnFS/LUZ1oKqpE/Y9Wx6me3uZrRp5HI6KKN9C713jQ
G6SOIBG5KlxSGfSacTkHu7Tm1NQSZ9rfYat6xYRsnh798oIoxPDx2G6t8w3DbJRUsa03X3cYIozG
YaDQVSc5nFBLK25+Lkkma5DZn/JtUglS6fndMcx22a2p+o+/YRkd5hpP9pVVbNxoT2OkRKUGIjJb
gOkJnFsxdZ2u8POZD7EgrYH37+n8hm7YO8BgJKr4CZ3/bat/21kU4hKuSbgwvDBKwxSbJRKsepOc
or5o/n2DXmsB65lqpbyUIpCMqsQIJfatZZqYmz9TneaQ2ajljh39xxgF0TZuhAaCsCLdS5k0Kero
f7xx1UqlBzBLBcW9qkMsvHdxPbgiRSFttEU76n0mbwN5i2PN41zxN697vmoktCTLljMIJ043fAg6
zITA16tVORfHJ7tSga3t0xcaq/m24w1ThqVAPKeSelVElJjwMrUyxscp4us4E3oOKmGRTzbCJwjl
t3EhgP6tTNv/vk0un3A0Sput2fsMu20Yzbt0rGro3K3rswKmCLhUeipVbgEGOY4lJ2TMYOTYi69A
eLocYoqYR5l4qpNNRtYrAbHSCnhTaWdfWc6FErC9f1YkhDE86Hqo41XmI2iekJ0TRdJ1ycUnXOZn
KNuDCTywaCLLaKOXEKaU5hcWsNh6o3+8fOESCzXIrOEa5PZ1N1SHpa/tLInIbp6Mwvf1Q9IS2TcM
mPNVr8W3i/m8SLGT2DlutsEyGVntpn3OloPdT+dDoAECWgyRfVWjCWfARc20WZRJOeHX8pWcCubj
FAfCZHsq1jt3lFGP9PEz7c05RPNsonumS9gBYC7pu+nnDZ3wXahcEubyve6oIVmMXV70+4PLsewX
3QnVQLjgSsbjX3ou9x4QBW9RkPMQN+fYQjgUrwZkuu9XQKe4Su8Fvhq5/y2PNdKMUAGYBhoJAU/R
jbp+nvfit7a3m4Qn6/LSVJr21PMlWkFFRDFRHy9RpuufJqxUr72dxWAB1Bc6MK1FMK1nIFGtMgVC
oZPljyQ4oqvb+Qb4YTfhUctWwMO+BUHt+HwLYBQ7N1+sHFRgt/hZvacZ1EIuwveAkUhT/HknEeRu
5uNWo1+ExtRwtzRKdXz/kpWAiuQjsAuA4/mLyK1deCUwXM9S0DpeR6qK0ZZ7n3o8Dw3D/wu9RWLx
TBXGldpPJupzY825CR9UUGPQQ+mwQNtr+MitA4iDkH5otvVtoN4aM3D62KFDzvVMdeOC0VqJtdVt
568krsA1ZzDzUa3iUAIbO/iquswSMl+jneaBmaP4x49dpob5WcVui5szB2hd93k4anQJg+EGEzM7
IoCd/cC42YcHdqUXqx/dTEi78hIzh83THrKJf+gFb46Pu4yvl/mzNzn3X0xV/lD0IZyovUtM1Ida
o/NkZBNws9aJGRDYPyU/19K/P/onOy5zh5yyC3ghBrIWfiKkJ6pgjfGPT21RNyi1dcJ7zgBWnSf5
8JznvzDB9wX8FnwdcSqEQd8Rgway865AErL/z1ezhjxh6Fnkor3BHA4Hwg+PYw4CSacm+yr8mBIK
Kl/fAsSqyE9ZJHDm5bWuUMsFEE7lrk37bt7vI/0pJgffR2gBX7ceNrVIfd8GqqWLx8Mxgcmy79/A
0OzxkdWFsOH2h0C6aiReHBz9OQJP6sEaJd3tlCDWbK6Wn8Tn9/HIcxs3AEQR5MzlTtybNIq4rm8N
I3Te37Yj86GJ0r9wJKFcOQpj1/5NGId/hsSvI2r5VmmxSQcKLTIab4w2Jnvdk50vc7a7Wp3otWQI
NAVW/vapfi1n997FYk1tbD2vImLyxXXlv2X5IGsSjQV5vue5rMNfDAwWqhaNFrJ2v2ZLSxJg8uj8
PujcEt53w7NnA6ZeLI8Jb2rUsIrCoBXU/cAzbO76GucLcmKUUkyt/eq8TWE0Yty5zKrn67bJ/pGh
RGE7nLP0Pc4hTu0Dxq2B2HwQ9YiaJiJ5I4bMEowqn++lbBkdcguVtDbf2UvPFw3BqjU4qer/KQON
pESLJVfYt0R1CSe7IJ6yBQgsEi5EFeUWKmopli0zpGxPwVJZP/lZexTp2tMzoHFr03NE2hCk1NQh
MBt1TWZy5ljuQn6uys0tMdYRsMueeQpES53RGNAHp8BOF3Kuw6vYDsDsEsJ/e5wFGZIQdb75Mgyv
5UpR8kR+NAiLlHkkZ8jlZIfOTkndf+v69gQpMx8o0dALXi6d8ZbVA0D3niSUL81V+kjC2sniccd1
zE1sR5iV0Pb/29tnXZL+qAKsbXeEg7NxdGxM/WpdkGyBSYNEKCMaUW+GDxWlxEgEs2rl2P+qgBGH
Ws5Up/YbshXhJlLdTA1xGQd2F9s5ArKxLu/XaYCOrQ4zjQP/JgbadN30XwvVwnyJ+pRGHjHqpRlO
7jhBmFBDQ+uq+M243+CNvxdRJSjheeIRoNcU6ZKeQAGUJAiE2ptNvVcevTfrRpoQFlOYeAsPi+cE
tt4+qEX7loiBc+5zQKx2hjexl5QbqhiTD/sxd1Z4P5dkIC3k2h09wBO+KTeE4tK2D/ZA2JN42VVB
+NjM7nm4NXYPVaZTCvkr0UXSozwM1L+TaJgjJHzSxBsi3FdBEGJLtZQw+QI+BVUpPkU5Q5GK+7/8
Rk6/O7F9qoZHX3CZ+2zLl85mg8aFF3jsi6akBUUjtIw0e85o3RqtrQGeOJ2yXi+tLEHOjDyAnVLg
8iNbPDD+RDeFSYE7BJD5ow2NBEGGTSoR1Q9pvEGZ0aCvux0hmGfmer1RDx466/mRzav3H6PAIASt
zSLdt5nRDWJZK+G4grlPrmuxa9N/26pXAK3QcMTgrcFLkT+9/pyUjTMQRxA0Z7ZjH8VRKO3EPRXd
kYLalpXeZuQsTd2QfBzVdeUcURwdYU/V6YgEFjDIRn54BKhClvUCZabin+7I1UPbz5QN7PjLQxtr
pSH2JZnCGDKjB80Rzj7J7nyLyMesmxdZFj0LbHjgtqRwULVYkReucnwKvUMPnQgE0ygVMvDzsOpg
Xei0L0iSQ42HuTcmbBprsEt1hQ0m6a2Yci1na0PomFD8LG04aa+3o9jkh9yzUS1Cp/LUOaUR6zRa
pbVmy+ykps3R2V3uA14JzbU5Ocui481I92v1eyYsfpDBLOyqBDEsO7P5Ha3xx3yQN/O9vQHbSkWY
0vurIgMnCaiyeDshVvKTcQVXRBwoBcQaBHT/yTEsDYTi9rnIk0C10MhGPJvffSw2WIEwTUUrltjy
1dOj5K36gq8E4v5Rgm5+fHAvglltNYakb3kTg+BmL/AFJhmkLSC698gUG76joRHiBV8FqUMZKgfF
KVXf+De+T08PuISdD47DXacsSKkjOzueXcOfDGd7XaIoTnqLE5GIdeDbpPR3ghae7KtCB0Uv4To7
9N3XGyiSn/rmtiruj6612OouDLTOqxTWiY/mCL41/z6l8E8BSl4VRPdT4OSG3eNVgAs1OE6MOtk3
tfq744jIsRIGzB0V84dEyretWXzXnS8gpXDQ+gMvJGrednucuy8F7wbxtBbeFL4QNv8+SMnFTBbl
G8F2WP1VifI1AkukRdC1tRGcuevZzRb32JSCa2cBgRZISxDJgAnnyp72HJxW3GVAjCPIJut209k4
+k5f5rC9HXKbwA+9cjI+F+U4iZB9tGEFjqK2hoL08eS+zdqXBh/nIBPFyxP/hPCENESMYftlx9Np
MX2inXmxVEENZmYlc6GK/GxEXEjVuCJ9kQVm9zkYYbHtyAcGaQUMw/9C9ShfBUaQXTSdYNrXH6yo
0eWAqKqbn2aLzIeTQeh7grnIxyvjOjwYT8o2u6fjoapL0h6Q2dbtuJorOS8mx088/x/OLadaw6oR
TWtocMhtLouyI0rJJI2w0Cgk8Pm9y6xIGGYtYt1DJjkZwlZN+DUiYhX+iivrSzr39anq73Jbzzgk
DjSK1BA7FBqaVCpsqMaOXRV8o+GHmMURFBVXKzuXRci2BFIiL+LquZX7hmzZebjTLgopMN0lYQGt
+Zb1BX7gh956GCQU0OHI1aj9pPZ4Y3GoERLx2LeK+fXeUL9zYktX7OknExRlIhB4A7QStlNHzLP/
Y258H9iHFeIpr4+iSAfB0tNGW2EOeRl+hMrKD7vLNzrcdoDH/AW7UiVV2nCgtDn9UA+D3lzzzl6J
sdyLo9JZtKTUaV7/wrTsrt0dQq4qgeCVKbySPmSjmY4gaZUtiQdwYb9aqgCARPtW4WU/4CtYxMch
1NWr63FUImS0GMD0s792LnwWGW6zRIB2o9HsWePs07DnFLzvvT4GSHbivqRktMj523kW8FBQuUZ5
tWFRmx7fAC5x0chDeJOiV4SP6FCwasp6+qDXfkRJh28MrP04NFFrMia7z8Bl/SoBeh0kTO4t40gR
g10doeN0+wudKw6Vc1p9oVJf7xnUtFm08ObTJhliv+4F3kWRKTysWXcKiFRTE6s/hjMyeu17R4re
+8sxHgQxkxVnSRyqb1mNE4JNzPbujlND3e3lNymuUkLTu6aNPyYfT/KbQOgArJaX44VL48eXUb1K
JLUBZq9OtOrlNvDNoB7w5vA/U1JCpzQhIXcGUqVnUdaCrgDCzeKY+0ArnTZS7mLyYcMqmp6lHL72
Sh3e+bp9D1X3lI+NEqQIBSzfYFeAJvlwt+Je1XjdX/ff56NMbpPFZijf2f7beLZ30JDmR0QJE7aC
8XwNJ3L5sO6bM4Zy/22PYJd0ojsHcupD8gy3sbjBE2/BSDSC5eLtFPsj1qASZSJN6z+qmdvoDsPU
VET2YDgUPYCYtZb0lb3fc3WU/yGu9SP880/vaAVym5L9SBmeyOGG1qQkHdLNVmuRJk0GSNtCB2g9
vpq6hF/oKzATemIS2ZmsaCa7HS0ggmJWDjJpk1GVFZ+aEJZaTPZaxDhZB4J8KZDWUyefPEE3KRf4
T/ffziLO5aGMutargtdVPrvOQiaieto5KdseEtlFSMop+eLqwDU6+ZpuIl9NE8kX7HN8uUO2PlAp
Qp4yF7OQeO9xV/o8hxuixaV+2HZt72oW0GmKxfw104sWuB2wy0R5sAUBGLd5mN4BlC5cyOc9Zepi
ur12UymRoea5s0Vyts+z/h2gw84LgkxIydyHl6renPEyqWtg2EhioxjAfzKt3pE28//fq6zmGLzL
gcA6fA/qYXJeCIxgRcXqDJtbCWE4M+DhSqii6N9bTLXZF2admped2Sb1oouk3/dV1xsSNQddrq3S
4tBnWhABYQ9HC/fbmsJbL+kfnQVjvtzTod5kpBzKwK1CsXVi7A/c928yEMvT6URQvH/b59ypOC6I
ebQehdhMoSp842dNOJWmghO75gIJiFaR6zz2Ydd5CKY+2T0F4D1uYjjvcupzlGPT5nLsfl08VoA3
3s3sYMD8OfNsy0dfGxdxAgNIzMmeppttxg03FZNKY2JNe8VV/rO6gnb1FI2MEMXTzk4zRNzUFhZR
q2zE7LeMoDMQvPZtVJg60DVnLUdFWRD2hgrFxZVAlpeBvL+Vz5TzCFdDaCck3XbnRlXwrCrDqyXv
iElnBkLH1OhxGC6Zw1BAvI23r4yivgV/04xDBb01ITBKN0tZXyMI2iLc8DLyQbB7FiBmmles7LS5
CGvKBvGkiTrLK/n8v/i10BOYDhNq0p6hwvfp+Z4DuHH5g9sME3fcu/cDEJp7RXL8Exr4hEwoXHvK
6zgjKNxIwKpPQTa90eF+2KKMbVmnfqv0PTD3Z3cbcyEjN9QtKoVR6Au0cKNunphfguG/rgx1UFT2
qOgyjBH1y/5vzNI4aBXfL8b+s3aRQvMEXoMYWldy18WRrqZiKhUJ17kgxvff0wXZBhJ5uhsNxnXq
Stn1fr9zg/EprcdSyITgM0bF4dLer7MlUuv6GU/CV385VJ1LFBr/eRhnONTvqJvmAAslsKYx4GPd
Ysfiw/nFfui2DFS2r61KGfbALASgPsUPJu1f6R0F1cHUAUthwK+Qf4mHHYXvRjCIGVQ2eFfpzB7e
IodcWoljKf+NsCMfQzJ1MytIvu8fzJg+NQPCa/XQ0IMZEmUI+4EcAj16+SNga+X6fJPLp0hjRYUs
ukd4zDKFWsZq7Jh5HeZR5F+gRoMQNWizU6XotO2uvD1+7LI9nV0iVrzEPtumoFT12qHELUFp6LVI
sFT+9YB/Gh7wTqIATKBIyT6q58s3Yf6jqbpWCpx7spqyADZLUvjG5z0JzJiALoam1uJSYGlbG2EZ
wSiZJq9YLpzhXzjEMyolKwndr0a+EJcRyb8p88cvwO9EGkKzLRPLlGV2Z6j73yU4WGkG61JYmaKI
CdMT2CwGk+/nR4MiKxZj88bT7oaesbPIk40h46/LM/scXeC7tGYfaB0SQc/iEkiWxmN5ghW6Ggoh
q8coPxBJ3dgj4ZhWSRUREpF3HY8fEsxcWlvzSeivYVrDf7CyJwKB99UkJUWf0nhml7EVAaPFSMa1
tdwDGluZLV/r7x6uhZm6ybXerJ0F4J6kMH3Cv8DzV/beIRzMIyMizSGTsevfXrV6ylxtIn2PYaKf
t0rKJH+TWxXwQ+L33sz78lBu8EWNv/EU8TkhMmFvIlf8LCOqG86vgbIj+gXYX2hsxHlVUjtXW3ys
j9SVHawsAR2HJSUz5Gy2GrHLaU3tVKAeQdGb9Hhw+IeWNAw/4rZ3guFXPjW9uDDaFXRCazJRcsZF
ZQ9pxGYq04XBnnJGxSQ6aXlrCbdgLIpV1ZtBsj/INBbonGXc6h+DganQzh5u+NOa51vQ7vxN8zEc
clzm3IPcc0QWa5MK5Vd+zTSKmZxVfYryEMBvk/slonW1kKRqpMdKHtZFD7u4KR8a0New3oDATX6l
hmTH82ZhuXkecKfhdXwEHtvNxS908nj8K1atgA40BvhKGP/s5kwSVJnASOjq6GnA2TS1BYMFOiGU
M9yDKDzCh58ZLPqeatUIDoyQ0YspuwsCWuVBCfUmNN9dAAmIFiw5m+H6KBs5aus6zu2ECbRr0Dqk
q78SK/I+W4SRG+XmAE/oKPcQeXtyOF1a/FE+2mB5XmhEwyzcbTNRPyxq0nvoCbEhtkOc4qSYLZc1
tlsmwoldGn9oxzQ+e1oyf/1T5rdDoIj6HKiqqQACpvd0wpQKoUOPFSXXUfJpDY5jHd1bX3QeaAeZ
xxifOvQvmgFpuJd+IfWV7u08Y+mx2+SoCc7212bPkpWQtcgl021HxwSxCRVeHFdV/MWJCqBb2HDf
E0U6xnxDePkLb8cvV0cLn03b5cYQ0M0lP55hf621ErvN29HCpSU2DXFQbfzvW38fITzMPM5+Tcq6
6NkyNqlfHiesNCNWZZC6JLBW6ulUD6TF7o1Pv0ZpY7p5ZleMhL1Xfcdki1QmsMV11d4NQ04ltVcm
qruGknzhTHsLqXSNSbqHhpnGkBtFpXi2QWrU/0VRLjmVNjP4WNaxMvKi7s/VFR6O8Q1Oov6Ac8WD
vHngLMdJ5AZAXcUcVBbbR+9DFdbqONPD0ymjpzsRiFYpttlHazj7i0jJnAmnPuwXH8U0YISzNZR5
ZGlI2RcAXOVekp8Z8REfjN4Ddaji+OG84090/lYpJgMsoqOd5fgcn84/zElbC52jEFBNB6fNSxL7
IMIZEu/X1Eg7LdoIH1koNXN78Y/kXM2AFlliRlZHRjx7/mqX1gtjFMQbJOIxDNiawPhxKs33jbS4
N1zIZmXwkktWdRNqvRMwBTRG/xtdZGNb+WxXgq26d4owNTSC0WNgUXxxt0285WzU17m6hK26RLg2
Wv6P2s5VGIPXzkTwiF63fTHK9Op+98kcro937VMHVaNTeAZFGVkH3SFAo96QfZ8MsqjPF3tGbwih
TnOx0agSDzGiOYiKx2ti+Zc3/CfMzHulDY3sAZW/NGSeTOd0JozFmWPy4/gQ8WnkN+vANu7z3n9x
YqO/K4a62XgDW086IdeBQPF7EpMxqOtJ3qqk540iP+Tdt546sMiOYsCjv2ehmswcGMI0dnkruEus
A7qXY3tmvGdiU5ZyyU+KW766OjxwNlGxawOlAcuiGs9NxXSRIxBqRpm7ajMPun0hS/8TgHIQRTiN
gvDJz62vSOlUL/hYwKmaB+EqCPotGTHjxtM8xGSdlsih6jaSQX1r2kH0kv31bAvIXyDPDX3R+uTD
vtv6W7ySnGEMWamJmDMve0uCsXkJrXxkVi96XcSv8TYhpTzclvaADYv8i6zrZA8Psa8KiS/2+r+s
sgpeQIygoSqXIBas2TDVoj/n4iwaZ+paU2M/NRd8KqBkatLZKNwjWnaFfm4m6Z1eV8dIJNck81UI
HsnVrCKLO2g/jx3pwtbA21UhmFeTN6m53eKeQ4VDwqyFZL50HZlA85SLpgQbLbV5qWWyFQQXY7IX
Q21HHQ3p+EMJwYyH+TWviIGErU2mE79Lr/qeLR1BSkbqDGHMjgwnnjWpawJ04tRgqOh4XuLnpERd
SVRGVuks17QCxpsWiRUmBDdioP81MPqcHJQsLx2ezfECovsNkty0GBSXOPyx6iziDCXp2ANMuFgI
ZLip9BoTm29Hsf2lFR4KyyCTOrZBD8F9iWRyk/+i+kdDiVIA6Ex7pP8q0IGNWhYyWNT/ZVVx5Ahs
fyF7km6ON0nksNWUuYPDLDElaabrReqx1H7n9J/YhTHRxQIWits1NW6a5nHffV6hvMpQAbWPZWPI
lc88v7miNViyL76tSnXfL7Eu6+xY3Ja7C+xL5QPng42IYj3QZlSFsbUxM8RHACmu7heMszNBlgtA
vJvuXFV+HDaov+sWHt2iAPk01K/kyobysJ8B7YkDFIpEfob4aK8VeSoYu4oLccNNiF93uJreaVNv
45Vuu+8vV7lQEpzAWZg1vAFsVxdgwtRLmnNPhiuxrL3CvEmDFTsVB9mIqpUkjD+cNFppBkzlM9MI
JHGRt8ISdIEXM/3cUa/75FZXAVSD50rtcRWZbqhwBwK71WLUnm0vMsI2XkD49glqzUy1u7lb1Och
JtLJ7n7TZa32U7JbyKHdoSgyyHqRG516FLzQUSGWfamoQSwghRm/xkyTSD1sF7f2IGiilTmI90LM
ye77wUX2Zewqru+BQBQfk6E2XD5ueOQl3Y0guc0TK9Ecs9QzrX7PMIyxpxA4fXeOO/qxirKv/ppD
IRY/4UJseJPjVFA+zjW0XhvSDv/OAHleYiJ+Lli3umjWJg9sHY8DsOVwinmiEjP8zDwUGd5mbm8b
G9xOoKbOVN2JlnsNufJZjVDUQx57Hp1MpRYMZuMfcZNP5o+Yt8MxQAoJFDkfuJIJeXEgu2xozZy1
ijyGpSsRamIcscYpNHOTz+lPqPHAh4/y7PyA1RZTxa+ugqdiyw8Qye2JCMO9rcsgasv2CgZQZwBl
1giFjZJgpsHsZ/IEhJ+MbuHagS6GKzycnib0p4R9g8EXdvm0N9R2hYdbkqc4at76A5ZGJrYK06wp
by3TlTcSXcDrx621WsCU0anuXq7WMAm0iC9l4yzw9XEUumlcSuh3Rer+ifsy/IXrIzCNJkMy83sR
q77bC2vEsWHAk/Hu8GqgugodY62sTm4xZSFr4ljQ3ivjv3TOvGIBc+fWMz4satBbWVuSMBT46UOD
ymJU30lG6tOVgAaDxUzHmRtlKcv9qawT3ayE+fiVkGi2uIvxGq+H1u2Dacbi3wgsVtE6hHzUq6FE
wARcHLofsiNpcv3/2H6ClNegmgJ4BW5gKPq4sGv4Kj7PwKF2Aw9VI825AZlgcr4ZMdrZE8Y+kWg8
F+P5NtuCsS3gp2SYVxwB3P0Zuh5Y4dCgaV65aqdnR7yqodmnkrdN9roRgMVW1JympW3EyAiKDRR9
U3qlhIl/zCFZOva+ryu9GPJnJTC74DYg3wV7sUUSawFvUSd+D62fch4OQjiwguLDEyg/Uw8UvkPq
/++ZX6oEFAInY7KCqLIxYSdyPL2cGd/ggwvCjqxmvWT90I+jyhCctwb6H8sXZI+3WUEWNSvjBMUg
2qEibjpzslnzArdbvL1WkJ4NiDIHS2Ru04zGBIB4cGXVtBvmVEqVoKN90SLC245IjA9Bq88JoeFi
1fXO2oXtCeJzGbZYOqb57uovprZ9YPkAhIAYObO5M9pQMoru2ICJcL7ISYZChSd2tRPwcQWkDmvr
J8YtDRVelTtH8QVjp0CiNLoIyF0y8UCvBF1tZjo3XolkOG6RyVVHSVp9xxmYSxoZDGscFAxsmrD0
q/5prTb+qUAffoGrGTariFdQ/VbJShkiX5XpLDdQvGuBqtAN8sTx7r2wVjcEpsABzd7jmUu3zOrm
ZoK4xkTTc1ugMnJSif0pJv1GcGPev14LsFaRPEZi0WegpNuKGWCIoKq1wGGuQX0IbAUUeNvWNkSK
cpTyock4Z+tymc7F4FOfR3Fg6W3m26/okbklslsUhRuf5WmgirxoqP8R0QlrvNkEJG4X296Ue5iw
IyI0P6fWkYDiDaaQETEi4UPdSYBSy++oKEbiz9tfXKP5joOYoy8uz4UYEtEAQdcFOwotU1JSSlo9
Y6GozMFwK4cCtAUkun5SmTE0L3rgBe3wVamsjRR15lpXKGvaFZaTFHKYGrpO7rgLk6oucugDmHm2
yrwAXVRVuNDYtny+x4GdsmRpusD5wEQ++P69pkwUGrDo1cPuSPzhECzru169HuEoXC5le0o0YXp5
ictRH7W47xN5wm6yh1zzXQZbEw1iIikf/BIHoxlSGE2fgfrQh0Vf5EI2ThqG6cYz5CmnDYNSjEVy
cDmEpHflpRVjmeufkvb0FljPh/B5617zmqPT+BAjouJZKGrpehIiHh94WpBw7UvAKS1WkSyZAmLq
qzbDPgfVccO+acRrFYryY5nifmTeTbRJ3sEa2VXfu7vEUXNVvlAZC99Luiazaq1jMZxTSqwaddoH
nwJSwccez04mPtUG8Uhyrv9JdL0SiJugLu83kbAEdtMWEqUl58NaS8LFb/oQAZU9RYTvnNDJ368G
OJlcMWuPU3V6qPLVOCZ/QAHKkLYp3ogwMhw9gGSXNGQe1vo4hM9vhqg3lP6/CVWBWFKC8+B5LANW
LNmVNqWEpskNKPm6Ocudey7eZs0AVjF+fKJ+IWzg7biF/tpguxVyNhGkl4An/4vS1zowrNCIN6Qs
xbYs0ccHqO7s+oq2zvPwsp+4O6+UZDKB2qjtVaAqAM3TcTYKzyv7hRRFdfUhcRqpzcT9Ib9y7QSz
SktLA0QpaADCD6Pb3CuQkJcSRRw+WA5LIz8yN7JnTbwzvt7ZnXJHt63sMDrIfy0cXsPSTPYAMUUO
Trx46fomPFL9DYFdNasH9WfE69tl5XkZzABYUb6HhIRa2ZqcmAc09YU0ALMVg+EpumR0IpkR3bv9
/7HsfnnW0y5V3o0XuCCdYqHvt6KlKdKbzohhDK3UHlNgncIyZh33cvI1ifveusXpnovLRlbbInqc
orc+hOCzKtdvbhqRJSDMUCno09BmkUitr68BJJhf6NSMNmW31mxYMz6F+Fzff01xdELH4AuIRpfm
fQ14ntt8sLznnbBstGob4ezWuwHuJfoTOuGTPi+NopG7ZHTw4F3wuHGEi4z//nAZRpomiZBgcMjU
f6/yDkQgNCtDnclo/Om3plQsb5Gz6ag/+WfX9NIys2jlPawg+FjDs4bueNJMmP9DA1vQ4zzhKPpE
kkr2T9l2V84WQTSqrZyp4Fhd6mAQOJh7C8wClr6s8tigcRcSKCGTF37a7CTuqPyohtThzmreIbIx
wSI7AKwDsYb3f24q3Rff7amb2WZ3G7Rsc0WPXCzPIG1yuVCEzgeGPXrvFi+jgZfR64wc6ZOJarCX
U7KLGKVRDgQ4S8kBfbi2nziW8oa/xbelhmPUToNOHz/sUFZuGolRQQeOPvQYBaMJ5G8qmZfvxF0D
CfOeqP6LPnDu5rA1gqOp/4nk67b+DXlRMjpa+s4nUlgf0Q2u8z4QUP9Dmkxre/GJXgrIQ13eBR+L
1yDUGgLjnKW1vLp+xE4ORfYA0hyVOjnN6k2OOeAnthKwkv1JvNhP7XX6Y64LauVjs36ioC4SRkA7
8YjiP3IeW70piMwTbIeBuEYh82DO2LQiYkQnMnpeLC4WOAwOdXgslndt49a5K+7pOfbR0u+ci0xP
4vKsJoRBLCPykrZIpmdeHOryepYFkSEKqMijY4wOlxGPlF6toJL2CBItJlEfDSIHNGLiODhYQ0pk
FJfdb0ABY+vhN8nGmxy9JNLhMvk9VsYbCd508pp0cC3oxuTxHt9oydW/BcsMXoFz+jT08EbhUwH/
30Fn6DrVZtXtxBFRd6E0YXdq8L9t0tQDiqkhsZTYTlnBaaINFzV3XQPzivWpna6ME4q1mu6sHq/z
w2b9fx+atOqIujSQsQ2W/iDvBgG3sGmQtvqYb8wcoetYfmWQGWhzu19YRiLatN3/6jYDjY9+RCoM
HBJQV3ekvu0rKWIX6V+/RusdlZZGyvKB3HzOI0SRNOQcRP4cprHFBa9wjBqQcoBZ3+f1snygjmsx
R4ykgjAE1mD2bv4Q3CEzA/CT/Kjv/Q6CDim4ApOhGUqxQc9q2PCJMkEdwk7l39iCKLOs+YxJwQjP
23uZNoCg776PabxRvHGHYTz+W8uO9WQvtgA7BQHkd0O5WljCNVJ/hax/nsMsPTTIOGcslzwP5r74
C+VvgD9tznFTPvTdA2zPw7vTxBt1+N442Bm4q6lH9xA6e6vIfOO48vY/YVChck/G2zA32c2prh4S
q2RTZsXSZcXGarHcfY5lhQnZugGeKdCwbwQ09mVBNocd9cN2iBvZ2fqmzIF4gVL3yjsiRTfDDbxI
gVx6d1V1M/Z2MIQaBxsaApa1+6hAEyBmEUuoy/vE9j+LKBtyqXsdm03yI5icQFL7Tvq/Lj0t5RpN
Qa7z3YzF5/eu7OducN4j2ydw5kiHXd6szs07CkaLBvKWMxAjX4+kiFscV0G05QHdeliGH4EWACiq
Yo1+YTyOEwJL79SAWjuAge3oZvPRcLjk/GuJu6hWkkUzYRo3lZvRwgJmKEjXsAstdLHuquibvjv9
V5IV8AQLApvNE1/0CbjuU+DXegNAZCY/qx5LpEFc+MzSOp55G+H8vz8qpU3r/SilG9hlOgFxONqz
JxiBUuF2aQyqXwf3KMePJUTkQYns+jrqeQTo11z435GWaRamaMaxveL/FIKklz1lOf9H9xko11x0
bqavVjvwbBU8CDynnM6apeFoxgX+j1DEgu5QTwcYJ64Dob7V02fAKXk0UZYdulfOEA/r6yo9hT+C
Kc68X4nMJtY7+iI7SAwWcGUY5uN60h5Z/dfktw//700Z/tw2nBJIRu9jwWpY0FVlF6ZyezDuF0wS
e5UQSHu2Ku1IgMEHgaTEHn7g+jIpVDi4v8on9MOgG9DxZYYUA1nURCxGHznZHYfa+wS9hF2Hoh8M
ejyh4kFnB8XE1+saGkrg1+8jrSo9zl2Fkx5lVlnOOewJRA4lhGFq+pJRPH1NeEhoEFBZpiUbiRgx
+lJm6NltCe3l/bpP3ogZDl7BmH3xKSjFds5sps5k6yDah3UfgU2FeVe8ZRDjea2luWCH01yi6aZS
Zu4gC48ZTKrxqePuOE26M6/2RGsK80PjAQQTQUOis8HDMScioX7RFD5oK9UA1nFe6FswU7ip4ZCd
4LPvpTtL7QBnWvG5/DwEq1KgLcAgS0Ok7lLxxK4eobEi8YsHnYD0a0SgGEZWZa3JlEJSCQm+Db6E
Lmu8TEukADdQUuHelKjOUd5h30Qew8U4Nexouz1ASV35+A2eBHs7HIK0eyNV9+vklQZFXaz16X0R
SvdIxPce7hJO3glpbsaRZ5pDWBlSLqz/9RFWVx+sirwdQJlXgXPIPyRBGv8DKzDZG7ZKzAX2g9sv
DX1+rOl5XuFA7j39HXF0F5Gk49W8xKixxIbBlcJstkwVvIg1L0mSz+pMn8y1AHDun7XVX6x7V/v6
z+81Dj1d5ifFW+xJPs/aCmxTlLjqEpVq2fXY0KuGeXo0Hq1okMkYcbz/xJkh1BJkuana3b9NEFL2
y4HnNd05BIy9N3j612CuzXmv1B32uzDB9qU5B4Yso3wTzhhNYw11DYGIZNM5aPlmV8SVInZqSHQd
oT2ZPg24jLz6p1SNuRCJV58+1LghvpZvW9YMvaLhg57AMKneQJex2sx9Qr902bY0X4l01WZt/LEI
ZzCvSeuyJz/eacEJ/MXrQItdKLzGCVAvJAJJfj8xPE7TfrnTIIrUCtD8Ehrh3RwGSTPR92PJ61Na
BpRnwSAsusFNjzAJCM0Xn3kva1NBCzi4wXJ33Tdr4Nh5lons4dnqovb9tmplD3Sx9lvU8GtMRmqQ
jlO4doJuyn8gdwaQtY6w3OsAkd1XddoYHpu53cJ9B6iGFRmeJp0kjVnWIdmzL3+nuJ+TR7EQnaMF
YSrebedvf8YmYFALxXzTJjr+Xhgtpg+uNphcv7bqMBOzAHI8jYpT7m8zzkDERxi57v2ZWNsf+U/2
xbKAoYTXij2KvZ3VpxMfy/2hXBT3o2ez4rWcPdX1HqL5tzLxZzMfWaGMgrpu1zpPhrUVOL1SBJO1
aIXKkO/6IPYyOcNGGQaNqvRxVLZ94G+T93VWotgtZ6G45fYybzwfQu3ICz6J87LKYVghqzPT8+i9
QBcpNmfIdA5al4sPw/xl7Z9Rljrdw+6Wm4+s4mIvZc7FYDTWjgubumeMxk/WOs2VN8i8qVjlnkik
gbazsuTlDTeC5SD785EF6smVe8c36LBNVJd+T/iPDuBvMEHb4Rvh/XCejumivKYnkVvdnGmIkO4q
Ll+iZhnd9s2HfKk3fZhhHal8wKIZOHda1vBEjPuGe8e+dkO9SzvhepTi4zQ7XvWVO2sAF99sM1Se
yjGWspesS5cCKg2dIFxEhSSfT2kvrkjZXgupOefqkcQpoytdu3MHS05s9CTnaRa7cX+y20QRoJPy
sSQGZoTEohHTldVZHxPl3HK/d33V4lSyqnj17d7Q6c86bXh9e7VLWfTjKH9re4scPam1Xk0KJnts
XM8Q4lNpoBLgSMNgPxgMaiLDO+1XWvdaldfomD1Me/6Il+P2RZaLMVt+4lOEAwj7OUmyL9YSUJyR
oVRwL0xzgmgh1CPOIL6ytQjnZv2jgnD9MNzyCcXy1GZRk+9m0doRK+8R7NMOxQ+ARgn5Q6MYk2yu
G7mPK91qD8hK2zZvvlSZ+qpzVmf7C/96XR9Rs/giQ5rtEz+sdInNE/ZbSEgslro2JyMT7jjdyyxc
VkG97RIXuYxLm4Z1d2wY998Y5XW/svZcMBvoMnG5Uaj6N+j5iNW2Zsftyz01fRujnz4PIWMCt2TR
rtMk7vkbCDB5cASWK0YG3V5emh9JW/8bgYH4rPwT8VbarMMRM9UY8yN0xAp2AijR8wkjZMUaUEKS
BUvxQZiQq2wSuKKvJzTsK+Bvf+316fh0W1Z1FXsVHzyRR0BPPHV9ulF0OIYTVmOX6CubNYDZnkED
b3cTQaaz/X8ooC7NBFNKNruDjeOxzkGs42bF206osGue0TdH/wo9WDRCTt2ZTz2Vqs8mNcdSeHr/
EJdIx1gove6S5KD+ytmIIJyVHHBvgpIZe2QFX/wM9KPPpmNjfgh747wsGTgKfVwhnvzpz8gjocwy
JtasgryP6IszDikEsf5LLbu/yeWiPup6b5hCkJ+Y2gpmVhJpgn4ZwqEY324csmikmvZCOge39Prk
BhTD/JWzxOb9Z9O38VNzCKR+RPsBKyR5DgSQ7efSmpO8SDIarD7gkpsB709OwJkw4E4i8QYY50ZZ
9d3b5Bez5LLJEghv8RqN+X8ffZ2btI02CstrO3MkhUT2MLsmop1cCGD6pFFeDexHVsFT54qeZ1vS
soF87c98nS9brpvKFIWvxT6jJao9tVC5tUrefX8MzYdiuwWBEeyShyaQq5c9bLvF4mhQDL+R8vai
rQfT5a/2I1zSEXjoGZI+Of5Fnw5Qd6Xu6c7TwKnh8tF0mX+rqWvP7lkltkGD5hw3a4LoLAVRuxb9
S5aGyms+QvYsppbBaPCb/7DSD06wgIfktKTOPtRezpmoglfFOJfKd8trNJ/3r3UbkCrkQbD/5ROn
VrzE0jmGMvzKuthIfMAyRpmFg930/fNWIhvkvThpGyLLHYKeH5BUOMxeG6JheT6v4v3QAdcg1YJK
kyvlNoMDLF2uZohfQQAoaPXvPHQXrNOnerIDHNMIIPvnsH+KWPayh8Y5rFUUKRnLbaO5Sg3XAQPs
isnqLTu7d308h2NUtXBDw8J88ULw6N8P5M53aUSXyHCNenwi/ULXPhfkAPVMYapuJbFPZmja6pKr
NZDlYexJA3Pumt3GLss2brb5LAEtNIbPe/018s6BfJpszMUloO9QbeWRgvEYERXy1iyH4VcpNb0F
WwrdloOhoF8MGfS7dSR4+W1MaGiToHQf3tdMAZdKVb8GM82QgGE9te7UJYnsOofbXj/y5XLfzsXG
BdP9W5U5Mi0CLqsuNyLVWiziminIUwPMxr/Qgxnkz64MDl+4xH82Ke5NniyQK84Uaa9Pw7K4mQw/
IvibhpUvwiXixnylU319Ve28KUYds+owtqI5VCvgj66buIWbnbiKFfLKxgHDr1DsI4HR7I4O1Bfa
lp1rGgt75WJbWDuotOYG55Od1PJXE0gXOtk+aDzraYSXrFBEwzm1X33Nia+trxVek5638D9VbFpn
lyhKBVk5g3reucrGlAHmLS2aqH+3VIaq2WpWDeRWwkCyzSWU/R/F1YtMP+ylz+BusnEsI/IbQ9+k
GYcajatfRLd/XG1LTbLmGtamzkzr3UvgkTYviCx40mY6hhn9XIjS8RQJkJTt3XkBBhz7LmmoD+OK
DFSEvACQt05aVWwGay8cMLZt/tXe87BdW4Q5Z3Vw+hYEj9hYNY8pYnADBTFuoHwMBQ2AWHr7kGMe
IIotSDk+P14a3FYMgg1O1dA0SZig4DzVpiznpFty9oH7ndFFH0RnGbVybj0neZ9IeQHlZpgtRGdD
zi7APspZMQosIodVJ2+1qsBoxm1l663AKzpoMHz8n/Tl1eQ2OIPyST6PtjkLmiYqKdpV9OnjZGtN
r6hL+CrRUZ3O+wyM1vnTLkkHafIp6pViHMu6+d/YTe4VAkbzzrlFfA6aKJyMyIJSof0rkQlkrtK7
EVRLo9TN/T7Fi0BFx8l34+mcafjxJdTIrYDJFCqU562BMDDvfQ2RJFGW4SoVf4cjEUb518FBT+Ta
FJuba7K7tJ+ZbZd0o78GHHtb4ByMnBgJWsT3zMVv0Rbx/kG4RkQ6/ja9l4PV6X/tkJNO9yIcYjNj
FNIIy2MEBIFTGGB5JlaTd7pbbBwznsDu83Zyv4XuBhcmwdByjPIgnZY/IpyXHYi54lnYsjmk9X1l
nm2BMtE8u8G8KSO8BJFw9dqIsIUxfhDvXZ1PViE+yMJdjjcpGee49TGimHyq5OtJqWcyKMGg476N
GnLxLXRvkQeWtHTgEGzzZIrPYONX4wdL5uBBzwSsxySbyT+g/MEsZeAZ9NGpBVGxOnWekk5ctTio
oXIrXl2RK4AaPO488UTUuBNPfgfqLMZc+JdL+4q3DsivVaTQ0bOtzwE8Oj6v3FCxbGlB39Y35cJf
NE5bqS5wytvlbhqYK3lLqE6hJxM7lq08RWKTGBYlFV8CVcaxfnjjKHjWPSGQkhr0N7SnGEgLLWNL
Ay8ogsQ7HHnZt8zOACqUgM8iOeFPRwgm3BWhCreoK1VRnewMveL+5xfZdkAZdVCKtrfBGRbjQqqf
3xT31x9Hr13ezdqLjhQe7URs/taAh7W2Qo2xTDSdmQj3/H4SpcRhWgrJrKmgYC6JYPjyWSQFowUn
PRdcX9FTf4Smu02u4Yz12pLu4BnUT/4ao9VKdZgr6IzewKts8861YbsnlrgHE55dGUUvSb8ryFcW
klf5qzQC+moxQQ3xMJ2GwmIfZRuh6fHFJLILL7wN0xIz7UtkrBkvJmqfY7eigSXKkv1Uh8jcrWnt
Z+I3SaGA9s2wuqvk+aabDLPl3RhLvWKDqauw3FZWuDmp9dm1MY/5ZqKzeEK+L/wHUwZQPpN61D/4
h8egqiXN/MoAfElgJUJPRdWfOiVFb4yURv/5T9UJbtlZCehEZhOPUO+FWgHmgI7SiFLFyvs+O9EO
XqZx+7ysX2/eB/F3pAqP2Zc5UR3Ke/Y5evVYezeMeQeeSgcae1/IVnJXeq3HarPl30obcscQ1VQm
elq79glllKFyTXqNLkfPIvktaQFWprObDwTjuQv8jCCaFuRzWScUYvycEJHw2Kw+3f+UYWEalSfv
5iLPrwOLOh18bAgyMuyNjuEs3kxYuwaJRxltommrQ69ufeZseSrdJ+TTpizqDCWMncapAxui7ncl
cvVtfp9xnUPQtHpKjHsEjldKouNXeIPtF/i1mfh6K2PB/OU8gPI4L7OIB3FvTJwMGKNLpe3UIOWe
Pd3X9Lx2DPAt7q6szH1u6Yhl0lyH5ms9S3FAP4/8kZ+iB/l+ija5V/Bgya2jVX/qxrd+PB04QW0K
/2Gh6EkSb2FAlVfsCdd/xxyQve5giwCB6+HvTsdL8QjmBHmCoZBoCFCA47APnazknYyCjkRNaN1l
igugB+cdDAnkOJEPhO6+zkCW5+zs6p63APAn1m0JSiS0We1kLFLEsIs4oaRwR8OZbrBBTEJyAgfU
GilhVKoxeQh5iX0gzxIaemzZ6b1ylFPtyUvYtTE9Z9M5qABNJrfaX/OZj4srucCfQ6lQE6NdClRn
pDVBFCL9wZXPfrOikXwtnv1f1WS6OOFjZl8NO4aRJkjlhUcomhd5NEn5vELshlH6HfxUAHq8BkJA
dh4pOb7+SmRNazW7kEh08IxFmMjWOAOlrhji7sQoVtSD1d954SezWJs4//nX12JImr44CZ3NTWoG
PPtiX58QY4rXLPUL/PltVSvRpMA10yuZ8J6nV92I7J4vFBiXKkJ+0LUWj+hUPxDX/W6YRKOfjPjP
SwOlDx7IX/nF9M7YHl4Ug+6v47hMkr6KoWULLQUX0W/tu/7td3itO09RCk3UCutwrDHQlE2XZwLz
TL3uIZPOurXVzWkLWDAsgTOCFfZXo/dUYA1kf685E6gd8stjYPQHWhzSg/i9HiCxCoClT4SxZKhv
WPJmsorAVM9Dr1xWuIih7wpoulpFHHQph2ZEEPW1TBKyLSJMKRNhWkWmhcGU972TdIeee2DpNKKr
5KHjBzFLaKCsGCWjPoklH1N1elmf2r/WoHuMoILUMu+eyabnRFWBjkhb+dUxKkQs4dSgSzXeLSUK
N0GEANiVXD7JJ/r2JCSVJsiovMnbhxc2vOyfhO49KTyd2qJ0c4HumC7e4hFwPTYk6yZ8R9vGTsAX
YKg9EL8WXi7yDs6e0U41mxKxJSPhY1XW2jx5BTpT57r2YrthI98ZOTtiSWdN4N/DaArOd+WOKlsp
zrXk6dQjUw1SYKEU3Ntjpti8dvTowsQNKxoSBsuaDY5hVQVRdGEiC/O2ChWbn+AOSQoSWDRZvq2/
b4PHncELpTgSP8WuNRiE+s6J6+ZF0YrGfeLEU78+ungjPc9Lkw2lo7S6ynHJPr/HJX2ctZfj+sS0
bdxEG9CgRpv0ak1LXvLyqMkdMGan1J4rCBjHFjEUf9XA/fCxWqDnv8T3G/UfFOPy7QVZ0V16RKnr
5PgCLj1hoeSif6bWCaO3s6duh2N/fGCRBK2JflO34+TzmvYvG9A7S/sImejz/b10ObS6fBzc60we
St6bPqgyw7m8oiVFJTZVDbOiilVVjN5fPhXbFpFL8SMdcFle3h8R0CbdIzxlfuVoN4uD0cHzpfd4
k6nbZ63XrRHourU+rtPwEauglDktkCvStqdfi626dYeQZ3cA3celzuL/SaaSl4PwPZ7XGryKXwQV
yepZz5UenI1J9W5u2bBwkof6zygLuAhn/DyA8jbFWnlKhuyF0jNcGvuSooaydXnZg2u3WUONmVk0
tjhZpik8UU5F0brDtfXK+qeGOCTamYA0OOAeyjgHsrKcRdTVzF/aWTPswkM3aapBrLwKcCjMjVlX
ROze8jt2cm5mC/WbaTZENllrtwdQ0/+Z9WE91d+I5fVOoS4FuaTKubYExRCehYHMU5Qb9fEdMHAP
2rIrDAOrOLVuJ1ntXigVBxGQc4nhhO6WgbrVavmec3OzI0mQoPEZ3jjzZl5wqADpZ4b6uDeL7wLP
FMBhpxfj3OqLjyJA9/2xVGsxF954nLEA0XSmtQD1yZmhQ2Q/F7EeTG0YS08T2URjKF+1BoDTEdgC
4xk41tkdooFOMO3UaYV+97VzNjIPcaTDGr2OiJpdUrzzHHiODlKS2x9MRfT82w7yBOqrpMlbIkSI
tASXpuX6y8z/q0AJx4DL6IEdmS261GJ1Ug/UMG0V+rN63lohtDIe32Tse3EAcJFxWK04jV1WSI51
c82retTpP1u4m/GP+mkvCB2zyrIfuTRfxbMQ73L5yNFzPUL26G2OzFmQoynlLEy4PObpJvX+L2hU
+q4sVGxZtf7NrppF6qD1jZ+rUahAYP2REadm100K0TaEz43STB9XzDxzQZeJ+WyyvHzPvEi/1ZQL
eIyP/kuRkn6La+4kBvQylyXGSy7XkVRwBVU+E2nCH6CuJF7EWWuf97O8FYen7NH1V0bCnGRD7Ses
ZXpiPNGZlbCYRTrI2LtJmfqRfIa5Jy+c6GH7KAKn/7XtAwDearE3ABf1rEYZ7LXDbpC6FxLc4CES
Iy/67dsxDiXQIBDauPLx7gYGDLn2W9clJ9/OSfxkkmyC4HiXWvRUr0wfUhPHgWWXZMQyEFGdpy1t
SnSMRDPhLhqYxn+IvVqZ1C8uQI7UYVEMGQZxhnSc7ES0n2Dtl1KOQkbIb1lj/9tlYyN3+YU6tbhM
+O2t95/9ovIftGK7lMoiOAS1m2zfruCaDmdQGMhqlHEY0bOBfi0tKSc8+J9zr9bYg5jtg1N96OGS
DYDdbzrkJdhcOsQChxdHaZZu9BtKf/j8JM/g6FLlJDCGor6ZK3aI2HnsuSa7gmEM1T/jOWeE3h/y
VgOpdjCL3moENV5Rwtq7VUx8nGTea2ATynFVSwqYaYaPtH68tBlvgchf+ZVv0kSY+zxfGr84NJHP
sk8RUQHhsAFm6L3ZAW05PCLrFEeB7cWeYPvhgOQo83dmMeRllbObUQGWg8pJFACjqC9l+CLV4fVO
7Uxoqaw2rd1pPfgv+zRN0M8Yk4S+0fyv/TIvH1ZS15je3CCPY5Um0AYVUXI40cevSmolsiWbglw8
PPUPxZrg8KZxxvzZZVg0kC7go2MMKv+QOz0dEhXIgkfp2lxQQZUoXr/80A7z+jsrnbrASpPHVRTk
t5GIrYOyA5cCYa2GhIw21N4IPba6nxQfv1/vpqlLohYKlUe9f9y8Na9DOj5uq+4su5/RE0nCY2Ek
nsrXqyBqNGBLNPX/nl1nhENFqs4Gf1Efa7N3UWYb3SHWm2nOhfA/T8XszGBbs8v8bli5MV+050ZK
/2yxFzpz+J21PPQiuFDdZBYbUR5GtIz8hoMe+q1WfcUGfWasfA/9xa+NmXC2LUGP78xb/tleBAPx
iDJywgZRa7dPIA72RkRHPEL/NNNyLBpJt6OEqb+I4felRIizaEf3rOlm7cIa+uON+kYObzUuA8Bp
p0nLxqrNih22mfNnPOdLB5r8MAK35fMil92SFYfylugtYkzXCt5koK7CPLiH8Fm9AR2kAXBULLZJ
LDsWIbe6w8niD1F/RoXhkCgBHTyQhTIFOfIevyTtZC1sdyERIvy94M0aRK9ze2isJTv2FEvvkQ3i
Mh2tLSZGYjg9k0VKFHa03Xo7hzf9AwV7/de5Z1ZLn9+buvOM5kvZ55c3sAZDiUyIIEaDc6yDtbRp
lvLgm4aYUKZ1gPhMKHgPwaj7si6MVF6v7Ov1FIEEjGW7dlNJojG+kXsBReEEx+ROZX/HJPZpm9mS
TvfBnqONggIxYKqe7KTjv84L1nGlL+rDDLZwqxYRl1mXZ9xYCDr9PGIF9uaygdPzewKl3b9HBMKu
rlHwLzptzzJFufGkrQHOOguL3fPh+Dh7kAquLbXODwFrP8k5gbkLS9BiF0N0ZPr1UUab9Dm3wKoO
gqUW5+p5xWcio2YUgG1KO/jDbARO8lhiY89umeJBFo7n+ToYOwe8sod+Uki03DrvxU23jP4+vTIa
uRQLEvmXWDRkpiIA4OSknqW2zUT1+/UY9c/6BwvNTi+CJIiBH24KoF5IIkQlxb9iESsIQwhJqIXC
V7dWlYVrsMk3n+l0LqNltBhXMqvuPIZw07xZGsFnFVKlcXAf2ZlXYnv6T5quGL5YRIMapSVv6TC2
eIPQ6++i/8RvJ81ywNwKdOd82L7Ry8KhpA6DSEeWyefYjrr2Kr/zPwCqjA2Jk3SJ7w6KlLR7TOjU
Tzkqp4RAr5oBCQZje0LPXWozIbAZMdIZbf6XTgyD7qEiKk4fS0MA5R+pkayp7feiSFX/AsL7CX7F
7h4ZzNRxd7UygmNPuJYRx0ip77j00KHXWai+FwLjambs0nYpNYtlz7lbj7lbCUOTL1nRTZLK4QKg
NLhZrxiKYZuTcdXn9C8yJYlRYfDel3SPLmwihqCjgRNRbtZufr7Vjcso3OG+VmTGGSH589/iS00b
OqTC9eXuFsdoS9uyRncAhSsCA94Qa4FLqiGc3hshk5JPZc0CgsphFVOou6DloiMDA9pw7RIIFQR7
Xq9vEQCJHwWGPtUw5r4MjZUY6DiXBfpfot268rMwcym9Wk80kkjZJv1yyjFJF1WT5kAqJbaKjrXa
/q1Tu2R/0wMneuFaypOOsMwqYjgmT9FiUTW5v8u9t8eKwxDi8CE5hiWliONLtWyD8OKBkC9CTfGg
ewx+VFd3NJf6oMQSTggUz1QLDhjvIoh+CJQghagpbqE/U1EpHLid/NINaxxiNs50E6gOIpytZ+CH
h9SGht84ufUJ0bhqJVNoopuXpgtvmeEOsmAcDGRjDplP8coSXXKLpr8pqpyu1gfkh8EkssiIMimI
zAXlYN3HH1NP5Rh0gasgxwiqQ15nbN1lVw7vRKpH3ajeyMy9NA48hVeKAN0YD9aDtdrtRN4k37lW
mehWjnDANV2afeZuhUOCpD8RQ72fDHKwjzZjZbUadbNc9Y9hkVvOEjmy4Vo312iFZTkOAEVRFZRJ
YB68vVOWUhUdEsXWArQlry2Fxy3GDP2xKfE0yZ83qecHwfwvT5Tz3oyvRn6R5zRzRgv7YTGKqifi
Puv+I6hhdN9h3l8DXzPsaCnEenxrg+S1deinuZN/msDaXP1DOEhOIqDIT2YwjG/P/FOOarmhaQ/r
NXH9gpmqspO8ZJ2n80X/9NinQ9Cl1bn/JjVN3wbux1Cfw+jrKwT8oWFEIqXfGrl9/9WOCPwMc8r3
/LL9jQnq6b04H1TUbsbBs2yV3saeA/gqwaIMpd/Kz84H9GbFW6dAQLtkIlp0pWMAC2JUE5Aa8Tu2
hSFERMUbeHziiEUGfyqqj6lfCuJNgYEru/NDFciH4GH0ZxiZCVn5JwXcWNJpMo/oQ/I5VQMWvy1y
bs+YR4xJvADwOzkKZv1lcLqM0YnSF8QTQdblRt7yp7XfSfcQ9lOC61PRM+NYho5dGYnxUqxN6Icy
MKj/+plTAvzvY4yAs3Oi7vhQgSp7TxzTKUG5myvlNo6F4Lkl1aVlqjdofZJyZ0OXDY+GMs0AxAnd
EkVu4KHtW6VMK0TRp5SK0jEI1BpXFF7YsGPWDgWTrBlElvoGX7txJKmk0NyvFosT3cnuIr/AwkLn
5jF/HoG/I06qoLjb5K04ceLws/YV2Vcc/d/AGWfmzrFqD/IpWhTWDjOJzUylamUsDybl8EdsAPph
1gbJQ3ToRvuVVNKMPMr/1dVomJu4s5wVcI1Pc6o+U7KGmfjRikFvg49nAS4rqol0+9AnZiDVN5k7
qlqiQoOVjJCX2cD9EM4hJYt9kWOFqmrnKdUYntD7+VM4PgIgO0P856y78amOkyt93xNp1+PEvdYa
d6dW1uTOXSkZjWhxz9Frw5rENZuB0yp8Q+KEn4N+qDbhR3MOl0a1XMFnW5bpSpB/J2kz1AT/He3l
KwGxThghJpSAWcFIYWNtKCpmhcQzmENJg9loY2phllD/1OLmdyKm5RJ4o1aYdRRSARYAHM43w5Am
ZIGdrJLSeK0qvRzJYPnEie+wO7zk3zPnh8UeaDqMVdJlTquAcaxU1wFZAJXoWWwVeP6FPgJ/u4MB
Jv1n/Ypw3zbCQtSu9Ij4Mcd1emLk34xNgmm/Ek7+l+QHDt/MiVicXFgmVQBaHHkzdtBYNy7HQTS5
wzJTo7YZSED98wl9B/gv2ORBh2dknDjmLKpcONNX9SQm7fz1B9WISWczw/eJVkC+YRJjWiC6/Po1
ilCTyUrFaw2fWBwfmyUUIdvYReu6LD4AeR7XIy4M53/rrIPEW4ex2PaIBZOSeYU5oz9hRd2dS/xj
019EkMA2HKHObDy+2da0vePAaZxQBQyoqa9cq42Kwq5hjCjAc4EDhtrVmzpfDE1doqL1/pSFWgS0
BBuOWgT2ZHVA4+Gu3KZNV/vyulLB4rFxOYDvnDmGLhIb1ekMM5mrenE6xTmF0EA5FtiPX2dJsDOz
3Ps5Ihy3yAXT+m0IzuzS9tM6ixYEowUj3vdRMzwi2c/2m0Bp4523QmEX6h23HCzG6HI5GwnWBnm2
b1wv4ts89/KHc8CYWN838hubRpw+K2ShMRKHsTyBsold6Hrty9xHTx64JRWVIPaoN0Okvl3v6FtU
neuLogfVAUUyHropCJmhfulxziWHNfcFxBLMN3t4SmU/SuUAiSPY97D3isnhogSeAScxbMLXbV4J
tfK94kiXXuLhMrfyPTgyqxqJ+wGjZR21SeqoV51/5DtIkYpufZBZGQtixAs/nGd5C68ApA8mbwxe
nGMY5KCAEgSgnRH4z8kBTaYE1AivzazPTG1glTyfyiKDmnTP0m8Nh51l4US09W795CqLLpL9zINo
Q7cOFGEypXYRLjsmZPRBeeNQg+/t96H1Z4loNEOJGTXUHMY4kzu5UhwploRO1sITCRjTK5hRBu2F
G6H+RJuuNEqkXGP3mFh0+2cnOwQi3Mi8TOzzwByl0L4Fr7VlOAkZ2plgIDfgDFNVSpj7pAgQxtsQ
GiL8//ZS4lV7zmNFscp/B8sDMrUHc8ISNyvFJfDVruKFN6E2DC6XDJyK9j+yg0MuHVXP/KZfDMWk
Y8LYfBfPkIrZVcAy6egXsuEqQgVDyz2ewVFwY4I19dhLYevtvGnMe7ZFcgrEpnZKbJf1SE10qBrN
DEcDfYaObREBGR5mYwlDap+XMZP9SUsSWYeofXKugGEl5kUw1PQbnnHcklXJ5XapGUpJtBJVlfJs
zQ8bDLAS/UP/EGYLSIKwvp9e9hIXp5Ogf26wR+LoUN2sDjDYrhsFchS7I6c0tOqzOsqnvx88u6kA
DZXLiZcoWNAGGRG6qXgchhocaRc+w63NThnPTWpVzsQSO08AUeUmwIhMnwQ6w+HJeNvqKiZAsUjd
txIadib1F2hLWr1CN7bBO4sEcj7Lv6wZBhbKx6DiCWSM7ZP8uvem602+FaUrHPHx/XJXwMcaGtQA
eSVynPBQ7gxix2IkuuaYLcOL4yGoY3nraJuVzd0StisV27dF/5tBBJxV0vAGxgF/zz58tne0mV3X
eIbdfBt2YE50jB5e7xCpdcEVBpU8q9uYvUGobvaWeAu4ZTbJjYf/zl31jKitF6aGvYG4VIPf3cyx
Upw7YaTXmv3O1ufS0cRvnEIC3E6TWGo+6XPM0h6ER8YoGQ5nOG0qXJgdTFFedgI0m8AFoWkHvPcE
QcfTwqmabk5wctc24yf8kskDuzBAphSCSs9Zpv543OLRbLSmkzjlhb2gKOw0OjWnf2lplQSG746v
xH9YCwVHMw8Pn1ouNn4hnPqFJuv/7GBe19Gh7FyUGjpaFoLPkAn2Fm6vGe8xeKsf6V0KnYr1n4rs
NwSoTWt9XQkGryTmwyT9ZsxaVrPs4HFrWCN1K4DKLH7PYX4yKPCpEro3kum5c/D8Ez5mqVL5AiZz
tysv6K8pqYbcYv939UXVE7p0lH5nDHLqwprfA+HCjAEMIoQDGaSK2Bmft1yAikOIRjcM/ni1Ug6h
dnuwCY2no0wpAb33lSad4Dkcm9Kxo1yvnw37j6L3sv8GIVgaCRUmVBuolqJwF0eJFdJ8P87F5LR1
lh1xGA7yBcMistCI9uN/9xTwZhgOwIJ6ixXhCOfo84qClTiSpI6yAlwB52ELpX1m3/DRniSDGBSv
UnbRByb7S7cXbk+zi8W7pMkpjXZgUCII2FLb1vEDDk28sG9GkrjLJiA5dpgK27aQcOF51BNgKhRw
C8x/EvGuN39O8jRSY7MWAN5k+apI94C/3hRIrSAUzyFAqIRrV8glYwlqLdvjkzkRKdqRG9JO+KM6
ZnZRN+QVTBfR9lruZ5yJbqhz1NYgmp53RS4E2nRuxcP+12zO6F1FCwX+aMYK2jsOyLtf4+Q0s/v2
cNbVsVhQ4fkR5HWZ6VanoX1bUObBDlZCdlIkW3gJeWCwVUKtK0FHXqBriFc6ezvQ9u40Si8skgyg
R/iXnpthCNaKZPEiGgant35wD7r0IY9nnKNOg3mezfKrWNMMc9A1l3hj3KqxTGv3JdVs1KPQom7g
UHdGeGp2ElfirrUdWOay4sT96GXJ2A2SoWBzYuihe0GGVIqmMj0qwMohm/XKgnbWZ3npVmqA0bjB
090ASfB5K+OGevIhtd51DW5Ltjs2fgRkKhG2qqJMlwgrloxFyKop7IhJhYP0or99NBHz2JgJrFOk
k6Ey5T6z6alOqcgQI8cHHOx9+CCsbwcRDMLCmJ8JTxXfMAIQTJlQz683khkqlMaxruDPRZdPaCP5
tLvmWzb5+t35XXIU9U4NA+PqUxakgSW+aV7Rgq5kwOqguvHEMIAOqrIC4osrONnjgJc41lrprajt
j/T+1bgCa6A9VV3/kaF6uy/KG8JJQj4R4xuu0Epn7u2T0Mcz4gQ1LYy1lOlYDUqX+tb1K1AqJKJq
SlRzrOzUwT9cDqvLQNioo1OpJGcNFIBPn1YOJBL0+wN1fcZ4gqQ+fmXHXFDTBbOJabMyjtF2eJC4
YJ+kq+qq60Z2b9YQ1YgtuLs2Z529pvSV8I+uU2NIdze/9W5iSyvfmzqQxva9Dijlq1AIfxzrejG6
2PJBD0l21g2Zjae4d3L6B9EocI6jKyyPns3PVMxkLK8vGzHc3TyERY5rSIvwzkEk5KmjtfSG7Ogs
XTQtTp8+ITPyOwnrr/ZxO/PgkjJjzogi98tGPYPTkaPjZj5Gt0BxVJACbQK4EEa3aky3aFWgsXvK
JrPEjgtBmDvz/FGTPnnmg0pbCYt8ufN7+WfqhYHkzAUlKzFA5wrLpywL/87W13//7b1BEa+uMREC
Pn7CBS8q5SG2XGV/fiHN+EtAYo6llt7m5K509m8Yp5Dro6no0J4zn3E1E48RrUkafI4ccIr8iBvX
Iyh9NzWayfNgG9cyBqoPk6Hi+UdIZj7s+3Vx2guo1UPnFXkOv1Ebt+U8FP7F/SQIdZfJOzwBwRMh
WXPsiikbRKonb4qGFmwST86RbU8JbCFIs9VLWCvkDC92ZTZnM7HCS6shp0LJcVxo/eqDXUXmyyQj
AOg2md/+sSDf1+GahDZ1lF90Hkd7P5rPkFCerYbhlWqsfe16ETTSWwgF/q6k/zc8UwNhdF/8Vq/m
i4me+Mz2Nq0tfLG47XESaAcK/g9s6Mk/iKiuHTX3bd6WZFuSxkkAeqJJc6q++hvy2WE4a8hAluTa
MRq6yoEmc7nUX9xYKiNJZaldAUQSD1Bt/Q/6OJyxqnEvCwXhfO7+rGSN+He+liD3jfz0Hf3z500H
G1mTS3lXBRaXFIaS96AO/W0qZZhqnsPooiOumV98afc5lpzxwBTjJOVxt/N6Wgbmq9FSmLlbQWIo
izgigXoUQQWdruWZ4UE/YbnVtFtNx8JpS261ss8zIyjGUTzWtVwPA9cfpNfgyH0lbEo4ATCmh/Qw
DNKg8NH5Wji5wV2720ACqnOMY4IZbpyqF8CTvA0FG0wlrx+eT6u9MtLL6ONQUkXhkQMqvuHdW6n5
wMpdwS9rk+Mz3a9sutCv2FEf2Q7iFqGP/BzVXcOnHLBn5K4rNZ+XyJlWy/PkYrf5UBcyUZ6YB3/C
dFz9CPs2e1eBcpf2esJwzP4bF5dwfTecg68c3WXw0yiAUsdTUgKuXOm73+s8JHGMfbeXuTZw3xqr
VnAmpbUMcSw+qgmwAE8n5+vtar69zFyCNCqDCqFGyTQtJdYOBkJqmUQXKjsKRX50F+HgoZ3S0RGt
cVRcGp6VQXaf9f948GWMiuc/LLKq2IEF/5kmLGI1Di2qBCR2svg2vRmB1vQV+HYQNU0iNg42WvZ5
nToW26dUeuRAgHxPTnYvcwke6g+sL6GPFi/G2YdpKoojXzZfohPG5ifL+/a5awkwYeyDwpeiilJs
9+ESwaPgbrZb7jMAGeBv4ccc0LDhDwTz7EAf0M2d7Yswjmj98Lhu4FAqijHp0cuukvw5wwUGBCKK
g71G/5XG/3yTaMVJEPdC44U9BX8/2JepXEO7qKDBNBpeC0jist8oY1Xrbr4Qa8CXXYct+zzvph6J
go2z9HF3A8xWNA25EtVz4weh6nVfEu+Y33X7v/wHxAl8yjBer3lcEqB6OBmtab6OKu6mV0g/rE2J
2KkdAByfp061uoXCupL+6X3iTWEtfpS9e+7F1gcy/btR5FavMHYKHJkNUHyhHTDUm5h5rreKQq4E
XZeQprNvPbgB3RPszngilKTkmROQE5zy0fJ9FirbzTEMgG/dU+oWA/qT373CTOSRP9s1zLnrgRRB
cKqFgffprL3XS9byAiWS3Xa3yG0ylrhICqQR3NWlB3GUEfdu2+nlqGf4p9r0w2FKsF8ledyQcGrz
bbtknwf3wL2ibGkPqLm7UpQOGx1uQJIWBFtpJaAbDvcDWW8NxRIzgbXXzqbGfv1wIoq9zBhSkYa0
h9qCpyqK0jZYh4WgCFAViiFeXzp6eF6iO1j06iCLALdBvnmszg2oLdpvRBn1lVhQoK6OyQzfJo3r
LKLHZbu5n9FWsl65+y2VlksGjU8BzlHP/e3rPvOApuWAoWZEkH8iIi+1ROQQu5EyWbnNzb3z3lVZ
vapG+FekETQEtR+7ryF+qjhbJU7FvZC9fUljIilF5Sc2CwFCYr/4oDMj9lec27ikgKzQ89aYUcmV
CMLnduPO/PyhaurEMOCInSlFQfS1hSYAjroSndaVMjlMT6+EV0hV+PxV6VRUO88YO/uAAKVGm7M0
fZAKM5CQk6gtpdvO7dTnslCXTmsfWdiXjCK0rxkZfo0OnaxqdetlDABxHchgfmJTD6g1uGhYSFrG
UoBU99r59jP2bjX24qezKlro8Fljog1uIqMtH6Mj5A+gJQHevFSlT+H4A6JyNDum3APn7wDl6nY3
jCzS0eMeSWo0LLj9HJDkb4sl0RStoq7CzHx7a1j2+W6Uwhd3ZXoqgHOP8TzDjoNAbkaHyVDrJEIn
7PKDubmlO1ruvtCCz3awgImc8LQuIQDRH3HjYZkoy2FeXGUtKwKfoPTTQsONzNKnGAhEIufs2sEE
Cou+H1bv5PfBiMYz0Po+FOe8GxPeH5R3bmfEQT3K2VIZkuFmv7yB8OWkhPmOR2TwXZ0ZTeuGMNF1
SS+v0SzupTO2/zBkq6+/QvwbfU7X345HFNH13P35+YF1LnzU0OljHaOcMZVWHw/o7LPqD8kW601p
mTR8WhPj4ClOeUI5qJF9yJnY61KxFNAAtwbJdQjLQriLcZRkwSFL8dPMwRR/dH63oqSH38g80o4D
98+pXe+f2txWwhvmFwSp+F43uHsifvoFVtK66b4FqweEhak6JFLs4bF85wQxTg3GV00eYoKtpxr7
0ZYGSPrfhkNBzpxotpitfB+SRcv9ikaZQo9URTkPAtrrFQXa4KZwpVFgVxcdkIlUSlwWqFabFTkf
IKtO2qKTzC4QlMrZSZrf7dlxYuDEuUKkwsxKXB16YPixUe410FDUklx2kYmAmagQGw/7KOKb5Vrt
/s43FzWvWP7meiuxGQzM2pjjujc1Tk4t23i+pFVU6YHhtDoLU+bYiWL1uyY4fRsKbpra9uz36GXK
lbHPvofYZ7q5tneFeVVeabNISU7WqROWV+iPBClpjC0bmL1us+UdQVItFQJeLco+Piy3sYEp5yXQ
UMXTIAIhq/cmByeYEyprYwlpWng1CNL79dECUgFo8snlJNhFdvDC3BJP2kTGoZMmIAGkx3Wd9l1k
XjSDpNDyfHKDyial9+u/r0BDRIxyt2vhY4xHk4FqofB6lmJo80BeCJRAqd9WJN3pPsk+TPUsoyFe
7OZ8sWGNDrYyDxaDWpxzHc13lhRapcSj+iIMf7903xwhiYquXxxWTuTx1EqF7ouaDvfPfVgyuxcI
oqxpA/ip1RSDxUsDsoCpo6ZaVD/J4Evp0+CGMb5/kCVRNUwLQTp/Qkb7XB1T2t0W4m450tQP2x/L
9w6Xa7d/84OonlNSGNnpixm+79slsXjX1MD5kmeYNbP04NetwEWMhWCcA3uU+1XWUrCSZ0vMz0di
SmSfPaLK3Qaejd+DRIoRDpW1a3JDY8GwUYMyHeytc3zc+I3oEX4i76l6MO8IKge2cvu8kvf/PPmM
HSX/LJuvqhxjrz/pPklFpPDHx7D9Af0pGebfRbruNKeI2HnIZRbbVyUJ78a0uB7RWa6+AUXkZCXu
eMpNEjAKYHrT8FgLYfEAbZ57r41w1SLZmEqlh3eamqVL5+PRqP8pHzmZSYIBGmpg+MidUFYjBYEy
OUTbxC/G4MSkJdVX1fNnPLg8M45iRyBTGYrZAGSqu2d8cy6DOw0Hsdaq617Yx7AhBatIr+B1M2HO
i1bof5Uai0IdR0jPPnKyryBLaz2W5BZbX1Aq/FYLwObFuUU0++ddwlz+ATGChf83knTrU8gdBwnG
gqkXFuVXnfyDu24J+KSDsL6/b+QqEn4FPTNgldrWT8TFrGIsRiOGwj0iJWBK2fTTAn+yuGWNUiDo
hkvW0AFw2WrZnM25YhUW6+pt+sjdQX2hPWaSI/Vkc1nX5Xy+45rxMwB2roQYY0LbcVSBHE/TyZqp
PSNvul3KHtYMHJZAlQduTwZuq7d0uWoU3+87ZDUVeXlb1OFza+BctAVe+cexxNLmAIysoMzNWlFd
nw3r6wNrRmay3lPHtz9EdGJE3Wk8CnBqFbIXcZtKcF3MKvy8sQpMQJVofPPQo+RpaMF/NW5CsRk9
eJ+JA5X+5CFKx+SxXY+XCfVNg8QMP8kP6EnPv38PSb1WHaPqKDEBp6UssCZxQSM6GuGqwkhy3z5H
TGMNRqcZ4ME2aor5xjk/DSBGoz2txOUllg5oKQMMl/Niifjw/GJgqfopDsOAxxO7Zy8w/zfo/Um8
3uKH4z31fZPpxsl/JRmvfUyMRIh3gwSfmslk58OM+LP01fnT/fY4QHe7MlBwksvtMi5jQQ66sQQ6
9lM9S2ZJikrOJeqsb3kvK/bnjpFauzB0KKQ8cl3J6XUU5hvc3uze1oII0O34TyjUEQGS/wiKSHWd
YlLLSY19YmzLNjytuMdPsdpmxng4zOLJrrmCqTt+XqIxLViCui2VjVRfVISmEGtETlaZbUEUVvoO
wUSeds3Gu4eRHdlPYvQPTgGWh5DUM40in0iqJ0EZIfLwEEpPbScuUj0tJg83TdDUYlOVVOEijVcI
8fXpVC4NLfYmRJxywBZwZO2dfA5TXWgHLag8D+C1d5rsTfDQv/iMIdaeo67Q5ESwEOtPlSWf/2RV
ZOiXS6gZhjppxUY8Blh7gd50zguTGVIjTG7uVIqk0O6vH5vtBe8K3tIOPri0vfU2XqSNWToUnHVE
WDNQhz5r9ThlaSFtjU1zBKsYErOdMH4qEqLJMzBVvkSi2xsS7MK9npWFRRKVFOd887MlMMOYswqy
2A8yDvBBUBww5nhi0YTbkZN+PsfOgEfTnQqwP6b86l8CMxZ/GcCetqw9URICZqTUceV4fxd84eNG
zi2wjpMn3GOnY0UKRogX7mE1pwplqKMF4eA1Fh0oZ5325u6xQmccIWti6iHa+44GO6VXdBx3CvmR
zsSLSSBBsiwW6L5ENyB8Vc0omeZphFBIsCOATG1QCeSv6saJcuBEvV15i1DWNxGYeW9E8AFILL3C
4lsnBhgSgwr5DJv7QhjAKh4Bsz4CwPS1SEITye8u2t/eMjmjWf8HvzPyYdVTFZ2oTn6JsIjJLQGS
nv86pMr1p93LMbywxwSO8+ZkdNBdYQFibe1h585H/Qd8B6U5BXIAzpuo60xpda4/4Qs1RcLv1IEV
fT0uD+jW9EypnT/Ja0gf8Nzswbl2i76LF25weciReTzZX1jtEon/dh6XzbX+6OuVwVNEqtFKsO/h
WR38K0BRAC/NxYiymA+n/Z3iOq1d4u9W2UQ1o5zoVba5WDg20RH4NomEwNr2aiEzXAsXHZBepuz6
Ckj/X1ooUSCUjgqmm61JAp/g6WH7W/gpNN2Fxu+HY2QzoXTmGEcyLuSK6PV8UYo6g6BiKsDXdCeP
W4Rifnfi2h2U6sb5RlYZiE/aQNJE9T3cXSpkgTIdAhC4vGHKXGsAIfVGi/HqDnnqrim5SCjKIQBh
Dp2PXqVVmXCxH0zYJ1EEoY0unxsKcd3nnPbIiHRRzhw6XSBGImfQefFQJ/kQ7L+fT0fl6Oo70v2J
cn8X5c87bJMvi9PZ01AhWOQxWvxQZrYDuH/b/92aXCShzgUN8q3NS6gq7Ml1pt6b+j5XUX0ci4Ls
d71I3cKZoa1nrhSBl9GgJ7rezi1kYG9nMVafhDNuavHAp+qN5cpFRv35tysCuOoD2FMfgEO3veQ9
IXfiPPMk4UqrbmIRQTvjFum1FrllrmmFoF1UUizSleiksa0Wipgry5GRUSPwP0GsnJFa64WT1Q29
oHbagnZine604XfP37QBi42fIx+/nrwvpFyx8Vq5RJDhdzshook7VInE3kLYqC76+d/UFZUQiSlj
fSwzYdmjilu9zglPUoWyPLUBpBh7+n0ECYME0nMl/mHfjp5+D7dwNDHR2GT3scQeq2eVbwlsC2Hq
/AJttHUunTwaJsDIB5plW0jTcnirWxOPCfpz4i2eMR3ltVCxArcCq5QNrIo/frtNv3k4uARxnXHI
n9gjcJX//jwnu6CYDuE9C8RacteO3PQ8WLEIR26JlD1ok928+R5Q+Yctv/tZNyKugQYDrGUzMLlm
b3x6YC1rZ/sMxyhyt/JDO69S2eQRd6rNOC9kcLA0Mq9KXY+mdd2dO31kbRrH+XAiWPK7OsK2N6fS
M0XuRsETKKAcNGOrEEwRgzciFPhDpe0JFfaOKQGoOokqTdqnbWQWDCrADnNuBr5StaJSNk1KE3gH
EeIN4eWNrG+eNtfvU/ogyD//NmGt0gkC9QHovCRDGcR0npZUBPwsSqkmc3kb6dbQBY4whS9hihVD
u7mwzr72oDN00lFWdmcZtxGWv06LbDhg249YvM+c4oLWxzQDh5s+jvlQ9/JD5EhxviNmuOzrDfFq
C552WEty0h5Db1FafIeZ38qZh2ehZjFr39yqQa5zOoSG9Hizeg1FaXfI28y2a2WCs21yOXMAqYKv
j4PF2Dhe174YwGycwX4PO9kpI353rArgEXgHpv9reJqqFzTYYFsE9IlqD80tNj+sf57v63zWqH5E
l3ScDlFO+vVcyhDKuV7QWZb5N6T+aTJO4+zKUbBRvgvjn1pO3IdA09Icp52xzo+hratTIoapRE1D
wu5EaafvIC0lULb5Y9MwQ1trH/Rt5NjsfObaXCR5X7O6JZrMGV9JfpkkPeOpPIH4JfwUnGfmV9xz
NNc23Dv91wEprIvot/2Jmi2GxfcB1NmJ2/J3CFccSo44SWHfiUOBY0Nxgf65u28dddg+2j33GPqq
NGGYHHhzRZAOR1IoJRTW738cmVxIrQ6tlzzyg1sUD9CXOfjXOp6l/+CMfC4tWuTylc5YlMTHfrCC
KHPWNvwIYOghM1x+b52A/vxZvOu2TLuKDo9faDa0XQhRoCnhrLwABYLlUeDX110bB16I+1CJ7VAB
eJ9hqZbcJwoicB1kjqXvlk9tQ+iJfhNLu8Gpk9p7VBmoF3bZ8bqXZxVMHmKaT8b7s4GVA+2CR+7N
OXPEdXk1RoTt+WxA9LrPzUDfK+qqCHz4Klz3ZQUkMo0t8bLtz4vR0YOHR/reENTNfamiYT/hwbMQ
gKz/dfPn0MucoGufSsGooV1WGF1qaUze4sLHgZhuckn8XXdVH00/4s4pZiC7KxOPnaxuRnUCCyp5
VI74UEWXdEtwqs6f7gEwB8gVgKvj9VTbdXOc99RFQxRRNDxFghgq+EhW/W/Bn0J8WnTgPpBu44d7
l+fFGzADKYuT7D1kCz7+wfauBGsYhKeFnfFz+9DrUK7yawgCblrgCs243GH3VunAS6FFuTFN00We
ZcpkJUVBeTRuax5XAjltiF8tOBZgDD0UfIVc6KkTKxtUP+etRZFvx7U4YtzcCNo8+3vzQl0UW8p5
0ImXTtBGWNoiyxrpOexOu/n4/zEcpe+KJEzn6HLHvbQycGVeQAijHGVtDQyrSx6uYz8CluZSEs8M
/EkVf+9vs8c2WLFwo26OpNfdsh43sqtTmpm0Iz8ffMcHwHM2ERo2ayV496pF1TXaa19Qykk2O3+C
18t5G9AcWLGelF52qO6OI+vGs1TNOQfJZ78L5oXE+1YaWj1xfQFFi1783hXn8n2vZkinFwYC9p9i
viLEizG5SlRFCkY2lwNjD/1E2E7K1o91QtMWi1xMWgcQx/+63r5g8EZSsAB5/8cfwnmTocZg7vjD
wbcv+0lc9K9mV4RvbNMp/lI+cRoQnUABq/moDD0FoKWIEQ8QOkFwGRNBVnOVwQF3lcLvqNGbLkhH
roMahMl+WIi1Iukz6lfAOtQDNCBqS6QWEEhm8SDXPF8WUpOsems9NfWeIU9r4s9Tp/Bh4Qbj58QY
04spotRR5HWB+gfXtvu6z11QnsycsO02kBp53QIOcd9+cnkaLg/wM1scf2wwpUH8ynqbpzvSaaQn
WS9uPg4Mq/1IGMYzrfgPFcjohgrx9lgoNTpBN9q1kzMjgxDxyl36rV3oN/W4Ee2fe6k9JvWhGDKG
FrLPvxg+LGSZLD5sSQKBCUhG/ypNyeVshGml5uYpld7uopfMoE8etxBFPC4wLHzp2iVOy5aF9kHk
9fxyJtKn3E2embnK1LvZyQ9l2BOAc+xXNLBXm+03Tisxd44d3v5zaAPAM3rc+k0MlJSKwqg1FMd1
x+2tErM4VuYPgcpPH8AjfnqO/f5VWNIYOk8aPNa/lAKc3gx6JQ91GLI0aFjQkuQrTL0gqGkU4mu/
VMDcmhwnI2UNfHqt2dOryx3QhVw7+zEXzDWSbx4mKJQfVxblqdmwsXhfyQkm9bepZNJQAzSvwDEa
JU8V+C1wlnxBObjNjFPj5M4H7LJiwuLi2SBG+EoQbsRQZJCnNpAzCtkcimL3kGdoT/dpJbfeTYhQ
1KCXKEsGtumnwZ7rbTUj6MYYu351p9Xzcf9cC3BX4K8g51rg076nIZjQRJcqi9J1tyMSusuHtxjZ
f85Wvi0jt3tMMkVBYMOuhvhBYS73/IZkHJpF13vimobzjMASQYKrqz9sOYQ+Vh2S/NtKuCP/XreT
S/ZlqfapVPqpt+BlMpZObrgEVPPT12CQCwsA78GCOzth4SAwvkHzTN4CDPD0YwkbrbDXwiisbhzX
/6crSAz5tUEdpW3G0WROpH+kgGWB6O1yVNp5tS1xfCkG30P82Jg70K3oZUbS7JDgHfT8N+V+SC3n
XLAVjDqbTyyYv1YhiQqxd82Db0ET7LnbKSMQcu7ALS5uJ7aqzF7Ev1NRFIr9q4hIP0VnD58NAO2o
ZLEqKnsZnedE66AvPZkGFrxaLP2qBbINpigwX9bJv8gDoqOOh8QsthG8ikEZ/Yi1adWqCfOZjmEl
9qDrBYe+gTO5bUo7v8wqDmeYn0TnB/KGt39zGl7hi3K4qFDjbZr2e442PsBdO1lfa/4hFNkY19/P
zfWFIlBRLMF8pB/l4XyNSlMP33RxpW2hiBf8tWom9bb5If46ths4QxlD2Fkitb1EaH1aSXqHeSu3
r1M/dtowVkvH7MOIbJYZC6zXbqxXr862eLQcEfkolY8QoMU2ejWvZ4JYMM9/BQ/1hhrihy/qFwcY
aiS/8YyHISqc8bresH5czvfzkLLqWQUMSpKaAAXbEUkOtELQbUwRzZdcc/XFaVZLA0/FD051+UUM
m5qJgp00zb0fZWAj7ocUin5zxS5chBnbxR19ddobIaPk9G2o8X3WAzU8rKPE/0fdTyvGUtN+DEK+
lpZDzzjw+uebzb6azncKs9h17TOIAU2/5uWXPzlQ4BmABNJ+SDi+/9sq9sK8ZUX5eikXxf5jmPwz
dxSJHemSh5uKg3Jf//qd1/QTM1eS9CybXUKidkoAXH6eogKFJ3BqoGxJwyMhu1aM7C7hQtgYViA7
q3HDRIhMFJNkdg+TUdyqyntp7ohsBJBd3j9UN5BNb5UryyQ6l0KlL8elMLOE4ONQU/96fUa4KTFf
k+wHB4PNtZ58YEWJNN+Fkdo4vVnHhOdgnmuJYtsNMoN15/hcqD9nfXBypXXmZIz4wABZSl8MDKFj
PZ2sS4J/M8tu3ZWyuy+fmf18IZxUNaDUmelwIrOfqfQWdThv92KfRPNnGqNNOmXeyDDADfyf/26g
RExXkX1E9113DmhyEvvfyrEimou89PsDM1sJfMAWwmej/jzOWX3zWW3t0Y6OrpKL6nOfEDtGkZzi
ifS6cjjotDyWkLEo0T9EiqMgzWHd8JLHil5hTsVaCACsJe0TpMrjXYhZhb06oXuv/oe5GahL727G
OKQRll6zlWMbtO/YscN28d6PtQNYbMaIcCI61eSf5wWZnoe7D70JqURVU4IOniMKH6sG+rqGTELD
eGQcCP9ryycTWBgqOUrwVyXTS83zUu/swsm+OZilPjOxzG3iQA77JU7k3/Sd7cu/DTPYUB7mviuh
DIphx3RVz5OurzNRgAzTD8JbV6t2bBnjmV74FLbqJh4qwvbb2lczN8Jkjapa6VlIMhUfGjiauRb7
yCvVS0vpUOpD/jt4fk2zuH4TVZmNZuOKGvLKxJSSpbvf7t3PBcGnu/F1UoHQS014KVEstME2Qa9A
ywn8YrJOKuzZ5LGQKbpAJMJijeNxPgqkM+NXYgr6/XYMg2wkoYzziY7/5R1NR7Qin8MOW2P7z5Uu
9gosGZYISlPVbeTYs05+moT3+eT40jmiRVMAtwTv4Wx/FNQVPit5zZv+GZkOHF9LIMP6rZZpQ27/
f6E1v02DPHXlTAjmTjWvt44oJWU57iTPXrZLZBP4D47STw8NqnnYnC6hYHXL9qrd1UKH+6jKlN8a
tlcHyRADiDuXfUr6czcyJ1abhQ0MSN7GOHDKTOQPvHR2GUS0FirlCSeC4w3dJZzLtPzb0lr4ftG0
NaAKjUfAf/FzYU9V+5duWQ8uaT6qVrMI/gqqcMVMCKr1J8ilDXl48j6Co6o85XoFZ0J845drzhlz
mAXvjPKEfR26wNM4pa1ow9fajBq6wsZd8GQZWFa5AQ1AxV0wrPRjcr6PJb4l+Yib5VGo/8sj6z5N
BZucnCcU326OhtpwLkLMpxfjyuvkXdNaxGWNSFfL7B+wF1KIuRoc/GkESO3lcKUs58fOB2Z8Oyli
ze7wmlTAOzrm9FWpi7Sbp6rW+lsA77aqnNu+e0LToa/76rmW9GAnXES9FNmDu8y+eZcRw7Ov4I4Y
mmdKPdvkSCku49LHLO8QaQCgPxBgqEbgy18UrK//tQL2NqlltJBeKP+ibJxrEsz/gm3nhmjp2nU5
e9R1g+PnjjQCY4VVYAXC98V97acIz0uu3Pk9Zy2AlBN8Fk5r5y5Xky856rUb4D1xdcNYNYz0vUeU
fM2aKwwMNywiqRBuCYSxMftEnme+P86gAtWSl4Ve7WxZAnf1aJLvLqhLrVEYj+HSsXl5kBN3EZDu
w2O9VmiAr5A1ox31amdibYOoTtD2hahmvUyxWv5MRKSjSf+ZN2wDyBng8WLEBnzMMxEgBd8e+CTQ
fWmuO1pPuMK/+wsI8ivx3PBIKEKXBGH3ajiy+y9vBDeb+XcKuqLXOhkLVOEiGZnKfGG5zlbMfu5d
lJJ3kAIpr82NXfKpTqsWOlaR5lVHb0jUwSE/jF2pPaqxo5P45oFIEwfJ66b3kvWCmJOHgNhPECRJ
MnYuzexXSCSmyi8b3Ofm3WszvHLKbg8HCn1igBy2+UAAn1h3p4OHGhI4U1Qq6uQRoOx2vrIGqOdq
yzn+4iy5vX/3V5ntD4+55VLH922ltRzx/m1yCI3e5ETh/jOSjUft3n1J/pF1b4BdHienepa6OrCt
1rGYf1Tvobfo0NiSqFm5lUT8ou88IMf2Z1QG+2uG1rQygRCmyMxP585/SPN8kUILqZDwCzU8IuOB
/QZ0xVqKeqK7zdeHrQEYqei2qBmi9EpUNi7StPoWO2Bhg2pXA6DhiBUx9e86qZbvi0GdnCAguAV5
3T4+DzpneujwuOVM8p1uiiDEjzyXvGjwQT7GF6W1bDjG2AxbbIqDHR0KrpiIsUsJs5WizVMSOChj
pIWldTLmsF9OsPinRPXhseTcqLPoKQnc9tLJunr+8W87ijJfGo8w/kPXwusxlUEFFEehDyA9vgz9
GYVuIZNsNFh/Jq7fRTRKkvGyp3SDW/7n8pOkPabMq6LC4782lY1XnmGShARW7hAej0mxNDcxhgvj
D5NGgSTppqCJq/WNQ29VWx+FQv+7bMNJwVdUe6qC5vxwRLPMpXaKnTuNpRBIr03BxRT4TXtKbPHt
c4EZPhwnEJno4ra7yqlaZllXhynRoj46wnAc72GonroufkHLecQMYLl0nc7vVvkzz2btvcs7QJrM
btZU2M5W85bg7cvBI17g9/6YpRBEWAuxPIVfcLzN3svXd6IyaF2iWXdyB6dwjceeYn2MOAqWmmcT
ZJK5Hjxk8egQnTVvdUS0JptyveQ1cM26wyVI+8KFHNaZ7UQIvP23R6e9SN1AuKkY9blg6w/lM6Io
+0INQ4X1iULGLC46Mc6FOHmlxRvkoK0JjuA/yRgpOZuL5KpHI8531doW34lrnOz4JLFDUw20cC41
UuUw0ddLp1SZZMxeqdJiA8DWS3E4VBp8BLXRuTwAjSMEzR/DTSNzoRkyv5004eEiCB04xbqxjtVh
hfE8XuESpIgbiW9UGokAk5rxTN96eQYY+AY22IGFWyVt9m0YzLs7t+K9VmESq1YkbX316u1ey1+h
E8gwKJqOAZ0VE6661gRutJJFbc+rYARySwu6ARPWrrcP8GV5nGiet2e4liKqYP4HXakww9q+3pmb
5GXFejyb1uoKMSVAQUetBOt+Nl/dKEy4JOutGW9CXg18gvoj6xnyRL2o07dCU+k5462usKZJgu4G
rkiE8CG0xGqkYSHFwXplrn09fB5y0qfjZ0V2GQVaevB0aqQmWTvoJYdARUSXRBqhzJw/iV12tJ9D
f25Vnm1pEN8MZ5THj9T+XlOFJeTGQbY5e1vhzv3MjKwGzUyoP5aKg1GmoXr8hKSgBUS0ToSiqj/g
XV2G5/oZgnWfg4D34nEtq7vJgTAN9nw1iHoVbEqL+zBjHimOs9Iz+LyzKBBjN++4VW0v+LamsZln
PnWQ6Zlo81cIV1t2luhUaK7GpVmImjh2EbCIzWjJ/NvdBi1DHmdKCobp5VIX7nrXkA/Ep7DsCcPk
WvB6vXSwZD0tR7KJf1a7hRl9Ch+zut76LRjJ6HcHRF+2b496mnL/BWW0w3Yb9KkqVZKOXxwDlSD2
iDm/87k1pvFWgBhK/omMJc+UjTxlhJW7m5Qq449zt0h19mXOl56fF/D9BW1Lw9C5b1l0IBpJmnIM
X1emdihZcSpHbAnx2LpBK3SKcy2yXyLfgRVkka7IYJZdfH8sxr8G8DKerH6GlhtzrjMI9IN/Hnv9
k4rD7wMSPvHz0d2ymv4PPQKWbTHn8lkShTJEGxzXPidnCwgrzCdWUvwCkW8aFTFVqqYlIpLq0zIT
mFub1gWWJWWJxXkt609463v/ZgBCVyBXSAzrxBw23aav4SVoXxL8CQD6j4fiPoP3aPIjGk31JyEa
fd18OJseAyQscPpDSYFNlLpHAhjkE1fdaGiL4z14F46ThtoTPwYAo8jk3Koo+18t7RDm4ExZpPXu
yNwrdIKXfYLDNXOu1bajpAy5hs3JJs4WHcJM2904nyDaccrHbtYI8mGDxWuC8IkVZdIzpDQJDkLi
8RN7mkchSAa/mzDSdyqfcXnX7lk/P6KaX+7fGdKVRGtfFLbwoz4vxgGiATYXhMpB9+BIUBgx78AM
vLcmvzLz2jBNQpYdhq3AZGO5H2ZxZwzkV6N3dMVdQxzVWqMx0qanwrAKJYdtp4zzmUptZYNcqYJW
XvAVYJmZw9ffDaiPQRWhHXmXAHK03e1EmXgxnbD0pae6xzPlLE378wPBUhTB3Dr/ddlzXTbzvTY0
wkkDNPv7FW066kg2qp4StOVMdWNjTenHcOOPMsYXfxQJ+cEEnWxuU/kdRodTDqHBQuGci62ukYRy
3mTacDRHD4uTNpHNOS+5ECBHrmJuXiIxa5v4vaXcbO6y29jxtY6WcqBZxFhd7ce2NfTBGjTweZSL
prZYkPSUpymUfZ1OHhOowyI8io8N16NhhQ77JIoqRnFoldKdRkRALfyFDhxyfyW2BGn1QfNlx2X9
tuK8BptAV2YU737TzawNPnC7ry1ESX9sxIvidLh5sE2YU+YET3wDjRNrapRm/AwHVPpR6MBz1nZt
+/43Dyog71EoW58oQxQ7I0z6uY0CwAX3nOC/wYe4yTLZXwnz0X9ek5RPRAaFqWzNRowc1P0MVpOE
ZE4R+oxXyogfNMuhq+cQo/+AL/6uR9zg7I6kbVSEbu+6Wp5YoZtrf2ubTRPuQaYs+vKWUrDcT4Nx
iWCt6xWo9mp7Hgx2tzs7/oYZaNQO530XjlnIcY3gevFif/s5enuYjzVpLHeYvax9ywZM/g9C5Djv
gIONo2udtD+K9xYT6gV1PVLgOECswtO9478sc5tPekwNtttS/frG+lm+GrshsYnp+JzzLca3m9th
fEYsBC76pCZN/0HJ5gKgQIdY0E9Pamwj7uSkRv2/85LIZXxHZb8iLTZgmL9v/lAgdXMXRo6dGjMh
BWTBAJUEb1UZimint3TjzJ25c/HiJLsmqTwNrbeFrHX1PsUlfo70K7IbBN/mbWrkYjvT8HT5euuB
XpaKxU4OdyDgSiAXPpRsCwKufNl/oEJ1Q8+SdEP5tWiexQP5eySFuRSfaO6aaFZbGtdpxMKhGqk2
0NHB2LBMOftH8FNVU0yr9bXOUnCPUkYjbMlQmJMtAdTq3o0EDJWHh1Msd9wpdtMrHpNlJkXqqN3x
yOLIKOzdI/fqaj5uH6+qg2p08nFmsXMFClsRmEewC57S3XzgXcXLZ8e1II3uLO+cvita9bFyth5Q
jUeknOed5feB54O/NzzpiEXK/KKLCetsIDdgTC7n9znf0bWMr4hD6HpM8MgaHt2UAXmn+Yxlno8E
a3Yvap7y50YqyoGKErq/+cnvukcjoecfPz1fIbmFFRvZmKi88u19RCTte7c5tpZs5UvMBxew27Bl
MDb+T3PF6B1KelGWoCNo6Zuvfi++Hf/DBE4gCW9KLJWmrYQ3CpMXFVbG18nuhiBbS2C22xjpyge6
fYRlM+N+UZLNtFN4uc/ttXUl8I1qf5bbZ4n9IHeh51jG5aVDuYkrMtR7I1VO/UKQUAg93/UaVVg8
aKy5LDpt8un8V0I0MAQZ1G/R65s/g4upaq7LhXFQZWVJI9828qysf8K077Vakne7XM5SZdvvO/tn
1ZJ4VeCbyy99wwC+Mz/y/8+gGZfX49B+mp/8C77iuYNc6RPzw2kH9Jzpmvq7i3Dhs++0nOdzXB6K
G5RnbZqNa7W1RBWN/3WdXF29UK0aWEpo7KQEpCOrR3u2Q6EuPx7DdPpR8r13vARi+bIDt4UPPfLq
MMSFcrTY+YFOo7VY+Iz/1++NHIM9CjBSnkK6d9i7UYZlXHa2E8C+m+xXNIFcVWFoyvv9tvqADoSO
1E9Z1KtnNw1i68qoPecdahQB0BjJjXECbn0kI8E0u0x0BkXD306xwYzmp+xvcFKiwI7hAPTh5j1j
Rxw1vl+aAgp7R0t51IHKGGozu3mpmDtJqI/AQoJJ3oGGFGxyGvEnuxc+0MclLBkAHHnnShtPCDYi
mkeBr3sL2+6swvvFjJy+mfRg+5jnUGjGT0DfLm69s1rzGAZ/Po6DVasdvNrvWd4QkOPTBBjK34AI
c4104IyV97lTbP9f1CuXsjN6WnmFzN7ZeO3LiJpUDHL1bCzpHTBe/9eYk3QjteJ4eTt24pxLGwQ2
mleQJs9T0bZo4FoAYR0TzG40d/sTpysauKzPZLcV696V7AzUWqjZqO2Hik3ef+xzY5xa9gQbZfNX
eyVqRKTEBD4Zka7+hvRJxR2RYWied2DO8aYCbyrEr4MY/jlJUBJd54h4ssRI9d4h01swK84Nj/no
+Kjc1DjQthzEG+RjjKbj+SZ1kdBjsyfNoB0i2O6nWOJ5tN6PQM/vxK+ks/sDazueyLcpX2IgFDbJ
RzaO/znTbrrNmA8XMslakZkpua/GvWmti9xJJcL+L3wy2k9YaC60o1d3Xz0pHJ9tSau/7VuKj8K9
Z0eIRs0or/8xANnJtxjj+Vb7BR0Ym9y2WOBca3SO+YoA3Q7U0H3Y6SvSrZbPoqkJ1W0yc/TxqLEl
JHM1abzWItT8u6ycnUijRgHvTenc76875RUjKVJ7osFa8/4YlG4+NcJE3RyBleGIfZr2VbvqGG+0
9jC7Duu4XF/buWpllSg1XHPMs6HKxtw5ev4JeADgnN3xZJlB6VQPxRM7xtC6FVqz/Z76zKh+qsrD
mPkw9Tghb4bD0kGdWw1E43bGuC+uDYM9afwvrE6IGwdaTD3RMwv2RFbG4/HLZd4TNlyniHtQPtZk
S3oZDs6gvgSCRkHviey+4uASqIqIBPEA+elfEpjoHLdwsgT8jxnOqOwSGx8AqtkAxVK2WdjN9hv1
27Z0DUVx4bGEfyN48tY8nuPFuw83qeBtEeELoiEnalrznWI1y2FAYPtb3Z7Cn2LEfZ0ViSw60ms7
BQseS+6N5ElVJh+BaQFhjfMCYJ1Vp8827LWwJdxrjrWXeQa08UQvO4EMjeSGa3R0V0HdUeuaNUgw
SXbUx1T3FKxMLBldR9Xl4VTMKHrX7mQVdysNP1b7XwQ7+M4cA8GtYGgzEjf2Vp1H3Q6fn43NhFoy
d17tpPfEMGKX4IMxG4z/4EdZ9RyvzLJJexsXh38+vEGHQCOa5tAoXYwRgYuwuj2knRiEwsdgFRmD
h2DeumhHAorlqkGaV8RCrsh2fY108Smu2oZJ5lJ8Ol81PxYUjqqBXEz383LsY09aqZaeLXIY7+R6
yYIMAjiI5f3Y5QV9C7AQZFw0sF6ulr1C9STllIDbeSaHLDx4vZ2MBrfOnxkftNbKcRUGQkacPuVe
3gYeWHsqmWlIv5FQ3AQOl9nD1/FhRNO1oDRO2ZFtBrNsKY8BMa3O0jFWRk5/Vrw2vlYsYs44j8Hi
Rkx2dMMxHQLvgBuBzmwVyzR3sRrviytvE6jEfOSB52gXKV+5b2W5kZQg/WbvhMXW5Qzc+3MWsBSv
tr1F55lfvp3yAw7vAac/MfaCWE6yBidrbz+7Mil58/DxSgOGBc0jMnSKAPsEXFK9PCWb6gOtEaCB
xCg6nHMC2kMDn0fTBrq/OyI5m7Pc8e1zkL32xWNlq7GgtHE6T5NhF8AuKFhvRyevRUqxpwQSCjj+
vqilpBgHpKkGQOzg8Ry3gfCOCEAJ3O66/gINA26X0bJCWh350QFbZmPaWekk1Rc97N6gIEqAYBCV
7iddsZBuLY8zxuUp57LqPa7WD+7279XDv6ngijHR8Nl2WwxGVXlxCcHgfEy70EW3uF/r3QCKGSD1
K6h2fQXFiHsTviUVlYbQX0rF1Tdv9ruj5LpUOgz4QcvTAGOejRXrEU3Ml5xnuXiDd1jFVfKi1Ofk
0bscRxsWLS87sj3/BHMAJD2GlAxAlVjOxrCItwqnRVllpHi36ax1H1sDBpbYzAy4MNU3V9KfLO+q
X+Mxof65cAfFbj4xrRkJrYyMIGsIO8KXzjbYpUWAVPUtFCad0L6f2dR8QWY7J137mIU3Cak7Q3rN
kcYxoqBEekjbkkUefGpwMjxbdhefmxVMWBvM0kR6YNp1YMWucYiWJj9KtrEcXjIO5HIlltzufF93
lw75IIf0HUtbdCLb3O3MgAH+cVaJBESDhQ0qsAXLw6NKil9lN6XPtVF2kCtVjf6QGjHbG3iqEWyy
lk/mQIlBaKkjP+GeTLB4prtuDGHNQc2/GD78E8FlstOhdnoM2mrKEmGuZPkFo4z1d5EJpqueYnpM
mPU7Rau/VielaZKD2tg6A7sw2YdoPF0ChL2CEE/XiSRhHDbRtrABrGj3LArKDC0l2ngJYVyH+g31
YWYdh7Kcwlzk7m457WgveGPyRXKBBS1lLbAmpqEgGwdoCk7nCNqXpuALYqGF+MpA+9vIFHHUOVOe
1IEK0nhN2/yj++E+ysZRlkPGQZ/ArvWs1L5lc95fsx8DAtyjfz4cPQV406bA7vvezkBAL9RRcJzG
EIW92rYrXA1w4PkEuwq8lg6/82vzo6s3mZw/MTj+ZbZoCNz3DZ3KFVVH4oD2qjY1e4ZRH3PStK2o
N6UPo5b7gukDlLf5scVoyaq9Znr/f8QzaIZpvE3ukwzHsB7jPdWyZG3Yb359J2teW/AgxKpQac2D
bHgzwU0iXAqJVwUWavPRCJVvxvyJqDd2cEbjP0c0ZVh16417+EDvJdXB9barjIvx6iHT/5JrK9HJ
g8BBKtYr9my9mPJ2tcaQobE4hUI4BJ7+BkL/5Rj4KP/Gr8iOFP5o+BQ+vE3VWo8gckepUNhgDj4I
zXZKYjPY6fSeyO+wLd9cAV8p6YwJ8PSqoG49PJuBYSwIw2BzMP3jeuzGZ5UzEsvSDh4CiuqqcYNp
OkeBmVtWrHXgVv340EsIC8+TW9T8v3IDNuh2V9QEZhpvzsodLzaagwsehKzaQ5I767QIya2zY+Et
9eStSu+JnDtiEBdTeCU/QLQPbKLQG3SI2Yc1NuCWNLNiq+TTxTRvwOesNkE9KOctu20s7LvSpvVd
IroLhWaNL2v0vUE0nM/f+It1O0EFK+tHFr4WUNLSAOhSSEccd09MnoZnptcqZNX36cUmLW50RITq
Ir8PmBm5IlZugyYeYZcULwBePBxPFIbqa0keUZjFMNQU/VLvRFyp0P3VzYAWJYJLvEypT7jS3oAM
Bv1thxwLZKRlnP7HFRXuCz6EJGsjyl75yzQKKuADO8xEtqpTwGYkX3kl86J9r6IXrGVO+jQq63kU
19qAgdRzVkqDkWp5Io3PjSBm31CsoVBO0txTFxyhn5gIhwk4+0BSEKrWCxwnlooC8MP0TGHcWGox
nb1LXyVJyG95mPSXvHrOgADUS8OD3U4iC+sYSCPeSwj5uW+EsEw7UMrk32WgQuw4seGCM8LL/EB4
1TMPNhmQTKUUBsFk7KoQjxAPZFPgxDv7sVf59qLn3xSmJx4laqN2M0JYuPd6vMfJROJ0t/uZHKLG
+6PcwXQ5KxAW/Frcz5GGHbnqZZCtteLJEsXk9RILZNonyHW/AN5vbSX7/vMtrtS86sRa32wZW3AB
HxnYmiR/6zm5MH79kS8icnkEHtnqrO0bj+bAU/7e+iNXl8sogDFS/FxbyC6Dy1oVt6lNDc21bmYz
MQwY8lxbofptYrq2IZR51CUveLg7x+xVdZt+Gkh2nu6tPSSfn0xoz5JWYuBrKao3X1wrE44aA6Vr
PDZ4xzWnNNp+dTDCNzkFOcwJLjVUAFG85wQI5Lo2lGpOpypDPjJ7kfY4vbDzQ1svg8K989iskVwu
b8a46X+fWcflja6t2sgT3aKhoFkYfJ/30IlNpkqONmc3+CauaPINCAMi9MizmQgRTQj3Ka7K+ls6
6IvWpGCfkBu1sWR+KoU5xuc2eMRX+XZaIlFt7FIuR7OWEsv+DlDEs1jbXBLIsOpnQj3+cYHyHdIE
PO2uh9EVJmF76r6AoarLIjyX6T/6HUbTQq0VJ2rfdg0SgvpVLDovI9xKfyy/zagFyy9JSywzwNGC
jzNCFzY82iQ6XFR7oJsHKEr17CKF3+NA8/fAYtBhTnLpnnQLsotr6MOezP1E1hD5Vuywaftc0u9d
kTr3l7BbhqznVlIn+Jq6qwdH6ezwcDm06QZHeimMhLqrXXL6LyUF85aaoqqiuRX2C0L05T9OPWzj
RD4YCboK0pTDjUQ5ykyIiZUev6MaBYBAvg2xoIRyEw2V2L2XiH2DV+chFrE6KHFlUeW2IvO3rryM
/kre/1eG7fNY06J3SYsHgTr0sbxGlWJQV++EvbUkpe6ejqyv/DfXHmOEUeTCpcQl9JDB3hszstIU
Q29aRUH8H9c+k9piDh7jc6rQKY3y28cocxCHONBQQxN2w2qDTQYNCBtCYL5bXfSuB9Ng31Lyrwyn
aY+O1IEe4T+IsheAMDqp7K5T27nOPiSKCfY7MRpxH54jLlRXGmLhX31q+v9m+V/RSwjiZOlJQqcw
rGD1Tk0L6DOtbdYqpU77gL4GGs6vhUsat+2Rbvbj7MtFu1pqPIS+FRQxKhHt+FiszJ0mSs0cIXV6
LoKTnxF1KHS/HzfR8NuCySPV33+T64YG7LFDJavLqTrbCGaH6nwJ05gKo5LIZoDDGfkm4u7/alAp
XBYOkjyiZiJVt+PWRfz4zdU/eiJjpzppOs4dprqTZsU7bjSkgrPGTI6np/e/4AvuPAPsjQH/0H7J
wwXnQiIzz42EWk3T9fujRwdqO7wab3NaZPU3wDiFUlq99kN97RsZY3kNe46aLadIF9s4HWPMIc8Q
1kzYqpCxFkxB2YIjuHkbKv1JOc7f6IdXYPA2wVG/i2vUZ63hEBCvj+wk5QtoKp/vA/6NrLmPah7Z
Zv3Gv1dGDndxtUm+gFg4my+MkBD4224OhRz22DhoJNrxwS+fnj5H5LQQnMFlhkZnpHQZ3+/XYqpn
WSmR2Un5IPs60LOIV6HKnJuUt0/AIEgfMhsgghnzhKkp6b8e5LQdjPVLA8h0ztgfOsJZLCj6gHq4
ecSuZc1KTWX2skG1RGr4DtBJn3OUbvjqGLDzw6XSN8Dh5gEI44OiromxjZqIOXOwiKbzuXq9WhZU
ofHU/4ZWEhjQp8i3YBqrFiSff75WpEi9shQoutK7INUY/fOIIjANkVYEMZCKPQFqOc/geka0B3kA
lxVydqUX2J38HHDJa7teun6aL3Wvcad/1UZwHLUN5tWf/vdgxQOVEomX9UZL+RHoO/s7suoWw4aA
dKSdD6Qk5bZaxgWPwwYS5ojQ5MKMD63ZHA8U15HBJ6xEstbyAxOa9Einexzbi273swz1+Aal8Sfz
bcy/vQCHh1kpMiTIdCAh5H45wSOLPuzW2i2LUubWMO7xH4E+zGen941F5mKmIHrZy1tbH1LXKMkN
22yd6ei+rDcU3dx8FITIAEwXASYAZaecGIFmve2fCq4qiXWEMVcX+SWR5xWnVIvkNLfYMNP1pn9/
Bak55H4ecdMXNWb2Kx3Busnh4ncqeZ9BHE9PDzlKRRX8k8EURroes+uxfgMSseg+2M8QU+fzAmlr
UbDy5E8a8lnoYM7wRE7i1WQbNj8YObPAjxZ5D+Lv/R1ueWGckgL/pCtUrlC7ifUKEbyihVr/m96N
AV26DnIIsBh2fONEclmv4gvOgVYtC3Bdz74+UIVKV2FOCfrjhCP+EQzibFSOYpSymfGWE8tXTWue
Y+6S+jeBbmdIw618aYbdrfNBuCQ2lKs3WBWzt77tX4daUzqsggwN6s/7Bwo2WX7Rn+H/wlGIli1o
7q/cy+/Ky1igAi1JtsElB52jD+HtLiXpt8iRKc8YlI20dp0yPlVNVc/KRKmWbwuJwaElUaYf121P
ibWFClbsbKHdVnf0OdBzXyxrRCK/gHlf2qYj0qhJC8D0WbrtPUROJdnXuMQwMOkMcHjQKs9Xxp/E
9W8y5bCno1wSd2+to6uXcxMJBQohhj0dAGLYHq6dU+5Lr1oic9B3Hi+qq5J+5JEB7v7yBPF65WDN
GCPEIS02gka+MSkdHOFbdOwTqOwe6kwaake2WVMZi33fKSgH+e3S3cQ9R2dI9B9bziXW4DQGokAz
GdWE1vdwCJ+qYnSh0yryBf60JiehhVzJraxUsD7EBFqK0qszgqkbg9J5mbMK3N/Rv4UgaHDRSKN6
G22Z9SVbAcQ3eF78upFy6bTXzPv7Ec+nfWV6+aMs3BQEDoDlQDbzDxUDJV7aFx/lk/tGTcDSsJMq
PaIc06EbxEXLJG6QMWfW2aRwKCB1IsSSl5UqWRSVSvWOtPVHwpTtnXdX5+ZBhwf4RFgrkZADdijc
PbSf3763ON0uHRERRF17e/u08Ab5VB94nmqwVxWxTrV5TSKehr/DqyrMcYwUhAgOaePGW8QJCfFc
i1KSyhT47upAOUtkUdHhu+Gq6ucjoRL9QT+GHtTbLKzTrwWGo2UPKBhcLRH2nOU96uUZLMR6+SFj
FpMG8DBP+IvcwiiS3E8cVyLiN+8TjYB6MnBZrKT1JjQjv62OfQeI7OCT+Y+6prY52YfS5NvO8EY1
pKIiA5k7VnEnckAwpY/Sn8w9UfrKR4C5Z9t91oW4yWlLXupevONWji9kympYs+uBMFVuZypxQghN
edeCzPTWlorPPhOb3P/ZuEQgwISWA2Pg0L6rHTtBRQ39a/Rb5Sq7C2rSrEPoKQALUeMXS3+799iR
x72NP9ZYld11/8lcAEKCN+N6soaZiW5V+VMq63Fr1COXKA8G5SONqjHaUFLaCNG+iB56xJExr/Kl
0xNjSu2stzt+zPRsGaweyXi+I7dhtBpMjy2jE/RBAjKzh0yIU+SXmtTX7dnUUZtQB6f38YQo/ZDx
PlCcqDe/BUZBWUCrTirjDq19CZpWF6jVrYdy5+GO9zRNY2JGCsNSXk8dou8tJjZINrq3RZizfcng
89SQilP9KDKOpXFgj6xfm+I3FYXz60cYuG6Vk5jNA1bQSFi+DPlsHzRKsWq1BeDPvKiY0Txn0XrG
2FNEFmv2qZRG/zziqDiRkQjMCffzbT6GAMHwtzqJEX9OSbcw5o5czBU+PnPApwfimKbKFeXIj2F7
HZUZmylQFgfmPPi7he3sAAtgFPW/VXoY3eCH85qxlWb1+cMpHxOnoJW1NAyZbs2TIe2GUdmkqxcr
sA/kS2Joou4sz5f3fkjb9SXbwP0cVk4CvyqLWGkRaGzgfYfC8iq1TjKA+W47bHbjVM1x5uuigDl9
Dn83HuxL2imCqAn5ibAuzYnPTOrEOxjhf8M/YSJ7D1HlRR3+PJimL2LLUr9mJ152JNofcJXAneef
QbiaNXOFfUZPiTeaQVzwfHk9KHxPy/SP3ZIMmFXyjoK/iheSCggxbnnUpxFWXlDJmpeystJI8sz2
4HrttECOJ9caPHTyiMRJdWBMFavFjodDT2Sb0FIs6ThcySUMWvkTtWVgL0u2SZUdRb49d56qyi2N
WNUmeRC3fQ2LIudSFhfHpJVj095nVddWOFrNQpiBGyfpeJyDAKr5i2LtmZ2ktnDSRd4GcB7Gzb6T
tRcAoZBzJZZkViLNPEl5EjldN9M8kQG9WEv3mk7zPTdu4oJCmh6y5Vk5EdX0J+r9q/PqKg8+X4b/
l0pAqWsAOtxewWs+kz2dcbZZz/u1OAu4xCFUls05BZb1r9Ahn0P8xDm2uHpdFc1PLjkMKXdJCsbM
cjaq5Y5hk+2F4IEBrbWFOli2ryobgaSVsWLLdOmNUH6LaKBJuJ9M9Td7eJprGfl593t56yM48G2a
3EX0vgJACIp96SeHaidZXRjW+gDD4NIHfLYVzBKzRIVTr1pGGvMXqX5KgQpoiFS8j2b5MxMpb0uX
zU481wGTvuW0jI0NV/iglppNSSzcxOV9XZRkm8RA+FhTxJF4s7ZSXmv9o+X5iASDiB1N8dfAmYAO
ah+24PXkvKZHRViVKzVopa/sv1MPmo0lJijqZm2AnHN+bPcBt7xmh7Eu0mIXL8dOrP2e2xawXUkv
7JoCQF5QkNyfvo6uus3M9W9n/1ngiz6429Wctarj0zE2V5x1Ceks6Kv4k3HdvpBY4H0K0uxNc0k4
s9589in/Wz9f8rfy0Xd6XwTVDm1W/QKbEsGcSF44Zj2l01mSYAtZUyWBoJOf1vMujS4B7htvW0oY
hgiepMjA9X9p1D86ENOSSrKHom3jDweLUJ3hSRhDFfeSYWvu2jiRTRct8lLSx2t53nW3jjh7cyBZ
iNJCYy/QkKINyl3ZNcM5KtPMw+P97OkRqZwZ9bzfcimVBZT2nqzAQTbhcygPrrm/OCpta7tD3Xxh
u7JGHG5yvQwPidAM68csUKeMFzOb057is/feoHy09mN7Ur59ZKwx1p4T1GV4Qgku2pjj4Jw7rO4g
HnI8m3zePMsWqZYaG2MuxHgTkyG7GhtBG4X+x/SEFCpLiVoxwn0bj3XMwDFnyV9L1OWXW+5VPLvM
T6bvQnAlGkNV17AvIVF/RYEJa5g7qhfLpYaoYg+fTpyHjan5A8MDitnEviNkIBf5Wq+1XydcMyHP
czXS1pz1+o1PywZM+zBwOeflDJsMcYr/IlC7L1KDSRCYpf+sYwuNeyqKVuk4qxCeV9wvFzFgh2uR
nVV6oU6iaDaT43imbIEAjd3muVg3S0U7i16zapVe7iCmBxMoB+SaCwTporVIMsEglc/kVwV4J5yj
YbWCEbPXZqQIqnSOmtJu3Bbs6ssaqjWxicqOrJo+wQfgZPDXdB/tWtlkBwObxNe+ZTJzjc/4+a/q
W2AFcEzrunrqgBEvbwaDhRyJrs0HanuQez52I1DslznVKNTyqqGOrEQrOJGq0nmJhiFqu+WFGLg+
NantSR76mVIF2wxAX9AlZv2fwg4OtUmcV83eGpFpE6I35XyodFhNztuiotJoKR8XKTFm3gKu0SPR
ywJCBg+8BxDd5YctDAKrrjZR9HNEZe/53V48zj9g2wkMv8epzs4t9Fo9W78PJ0V/EuatcNPJLc0T
MJjiQZjxJJd2p9hQ/1eBJDxJtCRJBrARmQz5mkXzUYiujfK+VqNSuUWJhhEgnijPVqtUxDkXanu6
FnlLZ4T40iHRaoWm2gnCHTIS0/WNlcTyTLvWPTp4MfzreoYBlacAhjlKJvcqyXJnqku5H7OK/4hs
IjHf43Iad7pJ6M1vxF4M/VtviKNrv0nW3A5JppvpJ/F8YUSrlKKTH6fIs1z7DSdJIXfVwDiov+61
gZ94gA47ZAJNlPxP7J4jy5wzM9HjVWzlQxekBwuvItbF9NbsCKMT3yYBikS9RXeH2FXyKgYs+6eq
11XdF5PHYZhdoMkscbkqDN+Pix1u76wTCS6Y444mycbreFRUTTzsdXFKGf5M2EeCAchzBYCAsSCq
t4YtWIBJ92kbWKS/AW+D09PXPBd7ee4QpHc+27tRcECMLM5dX1nAgW7kfjuXZEQHaALqA+M/Ox8V
CjkvxTTIQ3jLrGCDsRxdiJlyxf2OPMunBs+O6VN64zEelRjakjr3CmdbhxA4m0Gt3V2OlGrHdJaS
L9gB72YYSV/3L2vx8bOoru6f0pADDyORPRn/8zlFNr1IJMXDk+GQGnxarXENnXqVenwbXZubW4Nc
yB1af+3SAB/B8hoDVWw9KWWVoGiVfQb46PqXSNmY2W8j5AE59+STD6I/tDevInrPin0AFq7Dauoo
8TBmkWyHKoiUGulf/Vy5G+iOLPyci2poAl2fz+2E0USSQdqSgIdLiLsSU4HxvoR93C0qlTyHaGN9
Wn/F/U4VU9D7pt5C+a3+jgNTsKAHGbfxDD0wwtncUgXnrJbNxDVJ8UP4VHSJl1bk5AMUrSr74hPN
8v/s2fvSAhyKA+o/USBzcL8TyhgsEmFjJs+SGlo0eH0I3+9lY1MiP7vMgZODuvYA4gibP8xLZsnd
HQxihAjMsigMe1rTJR+anhAY2vXWj5801q59f/ML2V7U3OxkcwcSDfZKvUMn9u84nncFDi2BDJML
EX06S8H9s4E5npMNqMUNB86j1Cis71yoYzd6HrYBJCBUKnvvXXWjj0wukcgrQ57eOVTC5jUehet0
JH96WsfmgWT5Vk+A1UqS/1HSzivbI7NITtAYS7lFsGRk5JLcCxNSxWTzxgVBWKUz3kLpxf9u5932
JkJfL9huBf7BqaLPJ3pj67uE34RerPk8GUT0P30N7ym4qVS36MJWCXxATodAvX36lUYR5KmRiSZX
zhqHzQ6ntLe2Z1tq/2fRPRpdTiESNif3e3OVh5TZMrxHxL945+HlvatZ5xQz56UiNfvUOxQNSUx1
6+iQDiPd/TC0XQ9Y8XlSjoYDi5zafkz216+aKQ+MHu7PezwqDdK0dk+3SBMVWdiNK7pH1SkxVaaT
ydh6+kC8VjL1V8uauJSgaNmfbv2XlAVZt0SD88ZcSk0EXAjlyWcGYRs7pcr/xmSfx3PVn+Ttx7yH
p8D1IeZLwhmkYkPWCyab2TTrDy/dbpCDVp9NxvkQw3NVFxGPQ2avjJUZpOwHRp3WnYQjpsBCASmv
BhqLe4jaQgrWC9ze85hk/kB2onj5lJKLW0PCtb+octMYKGyg20PjeY9nFeNC/78T9+z6JoCICX4S
aNK75N7+hvmauLL48bA5dB4g4qJ0Kc0xs+b0pd8fL9tkZfJ0HZOFzHuuu+uIFOpx+EZnUJMASLuI
no7EPapjanx9rC4/lnoxJpnayUC8DUwbXvc47Q4NwITwJrw0iHCwsXYA0ICkKR00RLcXCGttCAJi
xoq9FfW0b7aKfMLMPmEqejXuPHnCCTLKFV7oGuVVFGPaPaqLryXkK2EJ17lmKP6L/HgO5NOBPvuu
/N6O/H6OSkFHqa+KoZLw4JOSZuLNoel+Zy8e2LGeJQD4PXYUt1OUxWUzZpBxwy2E4oLHNlsnS58e
SDeWlxpUSR6RSymMHGwEZr3kUVpb6QEd2KbZdzQ40pl+vUQYRUmhGEwG8FtLTXUdM3uFZLsAAY1B
Q+FVaVQ71eId5vXydOj8rdkFHwUhwcvcDgUTXRqn0TxBIqH7wDdP5ueyE6zlbHw6H8YP2hp3KKrW
tEbaLYvW90l6de24CjyUbTgl+r4jRuEIVw+LVBJy2dOInqhqB0dODjfJEySdKdr8TG+TG+IXzRfA
rsNr4GUE4mImLXBJScEwcXElK3DE1tvIP3z0/IifkLbR0oUq7yC4yCVwVW9TcZSscMyafurYuiTO
y80wYZuqPHwBF1t8zD/+5e5Fa+23oPyjKHknDD1GMXuxoCRTahsJgjNZ8hUivH+fjoziHGS5CQMb
Tw6ZbBFJ2T03eer7ljRIX4tCivmtub31O5ld9w61vXkInCtaL+NGW/AZbbQNmmEwoWGf8Jj6W0Zv
i5wLTToNC8utnyv4olr8exuOUt2Y80D3/2giUoGK3E/UBj0LDOTO3g5xxfx7zS1dk9LE3EdYW0lB
uPiZtbXiRBm6oqGttrnLEh5v2tqF0h5OpztG53OrEKRhlAGwQtMS3FMs2yl5uJ/3gksZV42KmFX/
WBsUycghM6upMufIUbtavKwc9S8Q822v1AMS1dPrN9FOfn006PYl9iHfU4hOEcylKZXYz63S1TR1
+/wf6gzZ0HiLW1Bz3bSQsLZgT6SBgYUEqMBvfja4pS4pQhZE2/nO6E4Ezk7RDwyq6lb6YjgM19g0
JgkGVFnYwoAjt17/k+AlvPOJ2U4//OAG0HNw3MEI+yVIe9TsYiBx+GqEF9i7PWLHu3eJRhlP2SD+
aBH2uUJf3odIylkyUdJA9c6aW+Bv+vWGu84a35OwRoqkWzAhUqtZCI2H996uqd0GWi9O0gdUgg9w
5jMV6xSRM6H352ex9i8tViH9GdMRj7XWO4yxrEPc0C9z+XWLQmcIcQlJUgw23H+CPDrZjnhS2p80
XV+dDinxGLTO1n3df+JDuNxRfbOptMEcLprwSU9e5rScjJVRaimq6yq5fnuAxzir4Z5DZhPYBB65
FoWBCmirAzMgfzbKrgYWWNw56uaqv/MEYHpE/4rP/pKHez66XqVk09Ev0pAC7krQVExaafB+qh3R
tqznNjWyn//V7rF4uuAr/SjQszpNph4te9QgCLyaU/vXiBwzK0CJL29O1Vp/ud/1yiAfhxLC9L2U
vlqbBQQnA7DDkRg/FTEXELlyAqn3zk9ByF3ftHsSpLCG0atyQS9nAClvJzilqAqVf5b/9Bt3pyJD
fhWe6dD2H9CdIRYD/GFrbHmwsptYmyiq80NBPZMT+DiZIJFq7V/HwGRwcedwQfbCKm441fuPdDDK
oaUL40AXKxdnd+/TkmV0wb6t5/2jFgVdqk8041zJ61cOpdGq7BokTEeMPPkHFzGVh9KnHXMruzV7
ke0z0i3TrJ+tlhytHkq2NfcS8zl44CLcGzRr5yWXfuOVxbe7BQErBDnaZgSxtkj2G4N9RMB0UBtY
U5XMGHjDwHBPIRb0RycghTNkONDOvokdAxDqqnRN5ixsbGFF3EeU3i7OhsqdQJ6dX5yAkaSwd3kJ
wCoZVXlWHCD4s8bA7ileJqHbNvMVAgXHAkctryHQSjH1UovIzALktZ1MU+Gri67B6jT4g4482ghg
H3Y5B1FeZic2jmq3wmojEAUXUuIYijqJgFlYnKJdvHdDSjp7bpVjyxCa3dm97rWBaGBs+gvfriww
0iOyiDjoU81zElrrzxLD3mxFIjEqIdlq9IJi0f44eCiTEKkAnrNaPGXXEMxqISjrXGz2LEcGRDad
lSq90QS6qtyZAktIJE0zDA9PD1TOlKjloI5kg13E833SomIWSE/VynQIIYN22bGXK/lckilUt0GC
haq6PmcDvcd1RbAhlFNjPFBs9qIjxfbBlBpt4fdCtfVW0FtIZZSAamIypeophqTBRml6zc2kVVeE
6Zsmc5DlSqCEIk34AqJBICVyJt8x4aq9D9/AjLodLBobOX5l4DK9wg8ztEmsUUSLBWYxIa0FPdmD
oPjtZCnuam/avdp0vr9uOOqQ9c7zfqXhHz6DLeNvQenTuxMVE8UmHRd71X1cYJOOnvpiQQ1ebeil
geXZA/gW81bG6B1ywzzaDTBTjA4E7RgEBk6iK7KH7rkkK1Kkw4sRm4rWXaPClLkiU49MY/xsk9AX
q+62uNFoi4RA9jRpYpCTIsa5i2W5Dj/Bo/UAaCFX1DyFJPpy8MZES5z7vHcmllCNvaqV76ivj7r3
kPIqclyIeRR8Iq+tHDxBnkHaHUhjjAXO3r3R4jDFCY1ztCsF1XCY2igxTvUh3KH361yHYbSTneQx
kcw91yStd1J+vtD8ZPKR7I7YCop0sOWSeF+AmbkQqhC74HJ0obq04q12dZLtNp5HVQouhywRgzBa
QIZ8huh1RIqlBeHmFQFzad0gXHTuIVf8TmgbiQ0P4DIuBEjMUm7qaHaWmc0mxY2qeYyHeV/j3rl+
g+ZGtlN85wH+hTdrLYGRylE4Tmm2ORzVnIlpt/uMmeumvr6n/+8B893YtQjeegc3nhhXAj7tCRex
uqhvSco/wX9Yra8I0htU/FaaVPJK3Iozwj7o2wybydJq1GZkSCo/yHPqhVjg8vz9w3+ehiRHyg8p
KI5Q+aIN6AlddbJ+NmssIjSiNzIFx9rxCZk8n9yA+G4xEhI+9vmRa6R2uAAXMF6IgDhWe4Wx2B/u
5BfFDEt/RRwHhvPwuZBxoCFAT2NI9kg0lqbnDR4y6PpK78lyhcnapus111gYlw2v6bAWencZCmlE
B5hKf7EIu7zWKP/e68xply2v7AKh/NGQVueElomQTrQEj68h1d6xxp1LQVafcIBXpQkCkeRkEgIs
Jk5jl2GKaySULQqj+hWEx+0sNtCH0JOspoS+9Iml4bjZ7gyo/o0K2w9XAQiajD6x56oTItj7epX6
AIxzMF/y6vL3/Np7KhJxvkHd/Sdzsq9Wl0HaYgZyXrIoNBLjtivlV1ta070BqnjxIg69d/bUJ3sz
vGOqFvq46BPH1i6ZqLZ1qu9/l8huP3JqMpffMd9BITQFgX0OVYxONw87q/pih06MyMeKAQS+MPgO
zMVzG0nXCcEF4g2FFFotmnNQFex4aCJsXSNQz2yZIy3vIKb3UDjFeDHC2KUvFP9CjZDnuBeFZ+R5
MgfioPzb5bAB1eL2I8WGTTbAr4uMi9wu5yYzcyZt9s+wzFpR7E2N5XGCD2ILwhd5YFLSYtmP+YdL
y8tPCVLpIJNdXzhpTRb3ooZtbU+ogAMkhMD0nDqQ/QUNcgBuI6npenbO6hPqYjNP+qppWhCQOFrx
ByxP4+VxN7f0s3JFvvS15W45wYuer25bnONgAofG98YiClA4TB/c7rFSbs6v9jEV4lvTdDjV/Vp9
N7UKccu06HLmdibY68u1gUn53+99b5TVhGyjN/5wAapt0mJgt84asW/6aBdsuL+ioFegQUps59M8
z+99bS1AHd/UxfJT7tVdyqqH5wkIHwSvaZ8p4NUbguXTwXH8QmjTEc7NBaQI21MAZqqihssWc9EP
azvjJSMFNLN+Yv6K2/v4ZH8rJ/+caRm6WZOZGD4sBteZ+EuCdwSOskXzqyN/Fywu3IZ/yNeyxJGp
IarBOyh4wexGTcyMY55vJ5S8wDGOY1Ou2caf93VlrJNrr87i0pl32n0F+8KgrTEHqs+UmoCLGfyt
rwPlos+VSYewHdFtNk35Ptq9mjXy/su2/le1izlaXU8XMftRuOsa1We+i5Pt2+OeTxelHWjj5yvU
k+x14XmXiCBsD7UBf2FU+r0A7JgAXwwt2hxs/OrlJE9wiYXM9wUhNWQe+Vrtr8uZSJQm6FgSr1cs
feOR5+kcI5lmu7ZOOn49mFhWNZGfL5Gw9/626OAPkUo1e4IQZ7l4HvI/RTj4Ji+aZra66JkPEbqc
Xh1J7D0myHhbN9Iz350MWCGKgZx4+uX+ap35zMghme2qDW6HQyEb3jf+VL+rsOUmuwpbMk+mDiga
g5bJF6XplK5JXmwRaLXvTfOOkN4OiLZaw/bS6Rayc/gMLmcwCUObJPu92qGWNWYZytSq98iD0AH+
CdEemQ4rad5WmYLbwxlAVT804PIlf0tIN7ln3rST2KXFdT7koHQdVTsW2+lcfr0GYl3LSyehEJLk
San/u+oC0wk8otqVzfpJ8gZBPFCPVdwHrtGIqDTIDPb1tGflnz7duRvE7rgoB4saMe/sl057cKiP
0CxAS022dB3AM/a7x8B33IAIESrdqnXPqBvmxKRYRBuQZSRQXImoIp4Z63SCtFk1qGOkLUljgPgC
H5iWA/3qP0JKjjy53btE56F1hBHLkIhAXAqb3Vz5zzhqWCZdRkFfRrhHB28nr3/tpvy8JitjtZ1Z
zTiR9pGnW6eyhbL9wfM3vD7nqTZQtTgzFRnMPVXyz7rL9TfgDQANJIMU6fLUAWNvgyUvcSEpYUm7
VGKQpamN9/JSAQIgyDk8KrdFxsbmoLnKcVHKQfkijwRDBFXnVHD5NtpAbzPrn86Or2NYJa8sw04t
KfKqUI4EQcMJM78IufgjCmBtSADUDCQp0nb3bq34A1SOBLGZSwBVylmly516FgnTHO1dYZhLKGSQ
X+4E96mx5ZZaEfEHGFeRxEMh+LOItxrFIfBtsfEyrRAVdg3oAGYGwcjhxhFc6ecE9wAOXBvCVaMD
P7tYQYrQsAn1r44H66pqQaS5+T/mFlyeekP1x74iVqHdrFguObJRoL+dYvsK/IIqcWxvafSt8RUX
eeHTkdGcWz3P89kiLX6rKoyQxa5JXUdB4DvlS5Fxv2Xj833OXQNy2ej66o78xXIaNTARzWgcUwt9
vPGPrtL1C9OkRAelWjBNqZ2NhFck2KuSaxbWTlQW7IM3kg1mMqxxqmCAIwy9Tga6K5serM6hlrJC
q4xV6lnmzsRGsXUYDrJOknyKZcTjGYKHr4KSyQmHjZuBfxinE4tYQeOePVHkaXn9OvucAg6Vkpv/
9+FLZ/d6hOZpoOaqqdxQvzik0iomVIzSnPC8jFSq8zwt/BHS2IADGJhliW9ZSB8JzB3JZrRvGYOC
5Nb8MpKBbHzEGrRIp6ttBKp21UFIAe0SdQd5/DybLGz2MqJ2TaqrMqP3lV2KswT1TspKXviinI/x
WA2bT6ziLwMHAQaQVaUP/3YiAUaszMQwBX7AKxzGXGNa1fs1n6KEa4va/daKDRc1rqFpEaHIxAPl
IuMVt6wUBbG3I2REGrtKrynpo7nVJVjQj5awGd5bppxxC2dE1BAvbRAqcmgTCPzWuFV5p0wGiiFI
DPftwKGusF/KkOiAhofYVAOTk3XF7g4lE+PkBuPsFI402II3BpFWcuZNlTyBwS7WMAXoDt1UKi1h
s8xlK84PixjG4/HwCRgYXGiHU6KzOtke4slFVvnDeZsZaFF3FRJTcjBUoaYWs0i6/SLjlKo+mlF5
8GxRpw4durvdGDWrkDUFv4vdue0b6LhK0UtYLeLOwey1u51ETjAINev6uKxT15+Ug3phk4+OaAM8
qvHcr/g5QPa/1ZV7LWvYW1E2f4RHgdba40XrngNh2soC91KIzimpkS2TCHOeXeHg0kAlFnDYv/em
BZH2h8EBQVVTH2jaBS6O5VZBdQXJIzsl4AhOVGTfK8fbRJuded68m7B5HMv2psNVN59SZrlcL0Sl
xq2fZBUu5FBb1Ou6225M/JBbVq68DREf2YRKldIj0dT32GOSm4Jn1Kvq6bh40/9DazcYLFx716rK
7Im/vjoLQtmz76xJfDZNum5Q959mjmyLERFQzUN64kFGmysZmelIinPLDvQ01Ta38TjIt7dPq0wR
Bfl55beOEw2K0Gt/wLvdW5ju5Tz3KnIrTic72ALdlEsHDthBf8zdq3ZMrm0zjPij1ACc4he/VqlG
2Pr7bG1ayU6ODFVnILg7GhLOo44QVeCnK7OMUqIMGsUzoyMeaA7FOrao75fQNsFXlt/ecsj/YYqR
RlvUtMK4h8gdopmkyDy306h2c6YxeFltEN+HcG/jaHkdllFdtckcKMHkFDGR5smLsuRYlq4s3H2c
yF0uqdC03USSb4O7GJeZH03E2P9rE1+/6xlhTJxkXC+UF1yarSllpcua5Emu4qN+DMqBNYm3W6sn
9PLnHKgMsVXj/W9mwcPUeRkPfDvF8DxBpGVOFitG9HqSVTbBTl6uwAkszx/blA6nUQelUyb99r2U
eISbm27TgA2m3EGMng1dFirbQlP8ww8YzVJ/0Vbt+0AMrfHmzZOR5Qkie1nKyri/PQ2G2V2vnMef
hczsLk/dm+m1rH2Za5XCtYl2pOrSlCAoL+W7V4Sa77ohYeCVt7rf0FIIOw/ZOgb/92TPH8UKX7CB
/4VIeJkMaI/tM6mjEg0345SmBPY5BMHnyGm9pGLOws+R+fWWtebiNqMSPt3CzWA4QGf3fg6tiEtA
Z7ImpMgololPGO6tqOCm2MyNUO/EWi9iC946Q0JrAxwFQekaIYQr4h05hTH3IyHFpC9NmXVAETKH
T8rRSym8bsqhLLViQFyRkpoudjL59e/w+zid/I95cvb3p1WC2ZgfLhCWYgq9MtGBkjMpsMeGsNtb
efF97/qw9vpJV4IM9qMDCIDGjPC1o/PadZoMYcH8Q7Em9snfeFNW4rmgCiZ6f6cHIoPC2suAVlpC
0ThyAkt+QXfyxmWpOG2NEP1pqncR0tYEyit0mc4ULOAKQGOFhcDMr6IjwalQho++j0Ga+oaVYDX+
ga/g+/KGdtRkHI8gG/4ECJSNPq05sFfp0vaT1DIKnNTyygO9XXPHOJZ5tvMi4LdoBoQP6TGmSKZA
dwG5dZ95SNsU8lKzgLBQePyXBySMmSuNuF6ax/oPg8tRm7VxTXIV1ox9myVLSROgCGnkE0yzb6Rj
/SVV+iqGbABLmAlFqTt764sCLdPlaSYukunLgr34T6wQSXlOlwnVB3jnLAecLslaOX/LrS3NeDjv
XGYlWB4bphfP3P5OEqkOw7nYebLVdpNZU7vI0vck+A4iRUS6N7x19BlI25H1gt+sL6Nvk0H2A8TJ
jAccxi2giZdoJLmo5PkY9lYMzCjrsOF9geenF0B67YcVYmXHhwJpJgf8xPF53ztoRJlGHmEx8e7z
OvxrG2PnfTXzZWf6a4QhQxCP7p26Q/reAzwtFIsY4tTZn41Fus3/okY50d8mepqtSow9Mt8Jg3z7
ZLD/l4Ijj+BdY4ySHiwRRQs4onnzxd/z7510n7Frc46D4SmHKDdEj5GQGaOqkjOk/WkG8fA0mkGE
yWfpheLH/aFDU3nga9zcOPt7H71pRIAIetVQQxvKhJJFwmU1JFNq9ZpGo9grGqZcAgr+XesIYmGw
kivz0wViKfCgY6oMRZmNALpyfkWsD8gdt9tYo9J39krNi2zGX7gX0nl9PcE/e1Q2NcdG0+vdKh0p
3ktkegr0ThAsK6Gk76t+9207j+SKYrWhNES62GsWBkRv9XSqt65Ao9wlM4kXJR9w21KYXBMmEaqx
0cUyHjsapMjPhfxioy6ja+Z+LgYzPR4j0Vp+AQv4YNQWV3NRH9tfEAMYMoYfPtabClZk1asB5E3Q
AkmiokUCFjlNA2nz26lJv29jwJRfIX7QCPNh92nGmFBlb5z/B+BBzeflW0f3ApWt3FtKtYbS5qb4
8DeWT9X+zuV3z93R6/UibYWAVw6ri5O0jPD9XTicxA9g/voJdc3X74u6vEU8Orn13vFiE0cLKPJP
O9eHR0LAKMBw/VXzj4ES+u8zPzeA5OvJujnLibpsLc7DFVDMPYv6PqDyP+Q1IHxxy4iqe8GJ8q9S
TTUBtn0sGSYoqjxj77qzlI8NmWCSprxadSkdzuLnbxfCYige8CqGXVZ77s21m4ffxprLhXTLAUK0
8wrmJOt3mxRAwaC66JVJcyanZIpwU/v2aR9cOFhAK0gjL7Yis9G/R/G8QUrfNNwvqFmQhu0gchJQ
JICl038lru6JemJR2pyTUQlp1knKetKl60xjIuSrC9ufVwodczdIjBCakF6Y8oF6DYqUk5XDUmtW
Fi0of2sV90qLVpPx4x29ir1eIEDG7P4PTob1QztKvbSt55c6jzaN0wGym6dHcYYLMDdpCwUqTDTw
lgp2w1VHIIA4pTaCZlsiFQMyQ1NMXgXrWHwpyVfIafdnWT2LYhENwSaHC5EmYZSFz+J94NO8AP+x
LS1I30qekxJmC1jQ9hs2lD0a/osAZQdHR9HcPqQQ+DlkPz8boAWIdp+vakwLGBEgpfEOp4uAK1yu
L+q0dc0XDY0sYDQ/ncAfAG1pnFM0fmJcR2Y5E3jJ37fKJRKH4QC1UoLj5np/OK6VUNxjNR+UDk89
r97aDag1qBRHFKaO0WVQmfQo7CokHCDrtN+ebCPaCepklJgsPK2o6E7nJ+1cervTGH2APilNyuql
rQbePH92eYa6kBGio6rUcpnYNOzpnn63ehMx4WK1t/lV9f3CjTfLof6TW4/5xXo9RoVgxqO56Q3V
QRGRPgG9Xbj8yjwYxByoDsg/UePryVyfdUrzLfYsD9RkgXfCxZeMwKtxmutZ5f2sEfYsWAeiKmwa
5H0gHGCqAa0X7oGU7mJvS9eTVlQZ1L9Y6KhP9IjE1ch1gUBtH+v/t30m5g9NFaunkuCCRVJQSmb8
qpikFDChOKQRlevWq5SdDifwwMjkZl1wrYlNxlpj6yNKuyuPQe4z4ayM6crBs0i47C2G6aQ+8ftp
cUGSaispQY7IsqQmHYuEBOUgj3rK1+8Lfuc515ktCGliK0Mi/Pgo0bzx9haMgP40kvMZxzrQw1YC
gFoasb6kCCR7yWQk3fteuPDAY7J59RtopmPJeJFQt8h4Gp1i0j/Eseu43avDKgKSTznQA3EwiF/n
VREFz93pDgLr6L7TSgXpeTDIBhGOeget2ae8n4dwUr98xst2BNuTvW5DiXTu2CRhsV8y+d10k8OE
Fn+KNKcOjCEntSqBlqIhZki8R/EZM0kWkTy5H/Xvu3L3OsOMmpuEMRvYUvsxNhTeDWNhBb+0kauW
PeKxlbZgJp85uusvAsMT8r93gYotyAzxnPCipPxmL1BbYIkkYzRm8MXC1SLChN5NcKEwoVC7IWlD
8NmZeStbakzdY94bDm/fXUvwozd4V9dSVesKErJj0WrIpZvHAAN4qP9GJs1PAV1hFtDsHvkOrPpU
etoBeZwmHV1zsRmqwbI2mwBVes/5QDJJUmU07qVyAvZVpmNNo1FPLs2v623U28QJ+51DKwbu+IPg
QQSMLkta5sWUi4XJDai5WI4wZWDjh3OuT6gKmIQhQ/VGXNxYMUPZYCduEhxBsUxnXlZypuU0FuTE
RiKSextDY1L4mUHvSpfU9PORBI6F4getTGH/YD0X9sJ7Lk7Lhdiu0mQOjECVOih5rjgEgv2jOYaS
UOmI9WFSlrNuvgiqM3E0ASqbM3GeJUzcHX2XYSe7ewoswMeXjEkvI0arJU3lyBwBvawzdy6Upn4i
Wg7s8xy92SiLXkzxkPgKQR/2WBOTskkrhAyb15Ts17/qdXwZyEO+tyvXqZZZyiKv4EAzpVuAEcIE
Ppq+58GsLFLrjxkQxSd3murxgcVgchu5iF44USTynlfdOpccGZl7AXb6EEZ9YmqpSyqG3X+Q7zm+
af3RXrH7xig0fIZRf5pkE20P9BgDgqcExFs7eFPfukrQan8S+gyG0ZhHb0B4TEtYzIF7kkX+PUPg
Xnt9NQpyV7kOScOZfJ+c/j8IQZwz7mIFvsuyU1DukRw0d8VRl+j0Luib5PNyTQqte0Ubq6ixUsbn
AkcSibNJzr4Mv+mtKLkLS7Qo4I+6FY7eY9PF6+6vNCD8rGD+K1WkYefk1wBq48kDMAfm9dZ/aEfV
geOdbTvwbgTBqSgTXADY6z83X3hB1G/AJVuis9exBlhh3HCYYYxyGhTqhWTF23pkvyKxzw2JwOQp
KeSQHA4Isu7SZWYGaPQiCmwT1fOLpURSF9mKlg2/Ef6MkfeOCfrD3XOLeuwKML9BH5uNgp6c+mSj
ftBVXYQXiFZpDqBFVVVLkNG1S4gCsNE0vKfy17+hkaPd8ST+e/P3vqpKMDAkcFLECe0XQtkjMlYs
FKginiVablAVyzICxIAsRBZy9Yc/nYrf+SuNaRfQhPFZ2XW043qyp1CRHI4V+LvmHYMW8wV4I6pJ
8MhExyz9iEpofVQ3kWXDZOmmxE9MBqgykZqwkVcIKVcrhj0ernX9H1aXNnlsMcdVSgDD1Att8r2n
ix7nk8wVCllhFMwtVZk6Y/Z5jsqFpJqOl3I/bxZfN+8LUaMm4f39anBF05Qek2PGfVBJAYa47z6O
2F4/5wtCXox019HLTLgsUQ3n0G87U/m2CyU1jNmLPvo1Cr7oneWcISvRFvhTcePV7d6wSIniRyBP
S1+3lxI8mJKFzGMmHDMs88R5T/dM8UP3R97SsfRQgto4VznYE+WsHZ0R9jdqrxIPMN7EhNKY2Kbj
40/3ox6kjkMeEDrP063VFn8g9Ipk9NPgyUp0KEj0p1vwUKA1Cu6pxGnlVBw8ZMKARYd6b9ytSiKM
I2YYDPQ9/adRXNl8NQ0r2jCxjmKKJf2TvjZkfmPPCxCNs4vuvwuQCVF8tcvYaHU7RjNORsvZsZLh
kjMsoevKLsp/7IwdC+wkYvqNtwZFTfJS2zZZDbVV5eRalK9Foy9d5NXxAQeH3mbA56UzinQIzLla
d+KDha3KxSHbmBecaXl21CA2A93i/rJjG8mXdowDIeAL2bneCBuMJu53BVbXudaSMtW3AflkUiRc
E9dC3/MLZuTb40SRhdPi1g3DglVoNcd0XmotQmqRWEO73bw9yFEjpF/yLYS37Yy9IWQ1UhdXy0hu
LNarjt/GDvvJskK/6CevCcGJGvz7hIxnnKJ0AQKWsIKU+qmJxxcCnXFOj7lJrS91nLbkOsB1oJmm
PDwyO9u4LlqmX22zxoYrnyHmgTJ+scIq3TgTD1P5LheddR9rNixdxJZjZ67PMYTLansivMv9tf12
wkKXmcExfo/RJ7ERH+Uo/CbpkLlJB4ZefmJi5CNsV/vYsxoH5+X4EKM1LoVPqTz8NL7oZKufFzfc
6jwzCEh0KbeSFtez1ZmaU8NiFBkXGI0p4P5+fb1MnLy9R2F6X0L8lNntjBYWqgzIn8USsigJ1lze
ncG/9CBbH4Z7lL9Lnw18UfUVW+Dua3iry1pfTGnWy7HICWsTMChRbRJtCmrjhIviqzgUZ22K3+FH
LUb1zXlAyxJtNtLoH+fgCxQDOOQrI/9cpY4AjiBBeYS0AyDRAL70p3eukjtK4vamDC739lRgLJr3
+yccIrrxJvetvbfV4SstxDy6MS57JgrnZlSFtQYx2M4qzhjr630A2IRc9CXlKceyXFh+18ae10wZ
y7fi5nxWfSj/1gyYjZ0vh7+5Z4GCgByv3yo9HdwsCzkw2rvusPwCkYCmFg7wtUyElUjRFxGSENgR
KS39akhIHAPwW4jQmTB7c5pb7bMaSugrKnXm5mdYh8mLWYCcW+Tfeug5LkGY2S6HiyD5hQ8I00oG
NkdVXqySS7BPBXNOB5+m4Chr5KGNdlowafMA8y9PIWtqemAZM3Mz8QgqEfDnPWax3CPROVSlqtR6
4dlAtPpbxISFgRuvU4kohh9Ug9A72mawgsBg+sXQwvAT7GwC8xe+yL69lgueHm+Dejpr9p3n4jwh
JZA55sfVb8CP3RT+svUmEUFwAPziRatjiQ1GAvHfXg+NQw+z1a7PdBWixHmIqEUp26qKHXVcFJyW
z2fObwgVCcA9j/EVQKz5OrACJo/edBQGNwzIqzWmYBfPSEitpPWm8KseuCZB79WmAIkXHEZBoLTm
RKwBv1cSvpoz4Qbn6SUm7r5ep8U2oA91KGqbl/2ADoxI+xI2j4Erx/AQHfLuq38U9sGiTppv7Bnr
IoajxXVzYdpHcBwFqGE+BY8HOBJpb0WZZDN7NVCMaBeEFUEfIvx3jljXzI/JLCApADReE3urGyC3
qPXvdtOhojinp3dstGXdbnVJoAJVyjMVh4dgjR41OH0UAo6BsyXVp2AY9pxJLizInH8q587AaX2x
7fWF5YgiTYV5Qspd3PP/Kb7F2ZN8kqSyDv0gWVsE+BUSR9MYvVKhg3BhxfnsTVEbF2naMU7eOad0
3NHnI7LB/wcQLQWi792rY3aJJGznuq9od6H+sR9bcLpf6pdGsUBDD4PXRjtJjfZiLTfjFGJKWLyO
BiOyFIo6NyS8lv1f0xroCRlsKeu9U1i9O24NflNU9Laq49jmxSM9E6kgk+TcI6Jv9R/kHja3iaTZ
0pHpGf7YxVOb6PLi1ugxD7FmULHLAKEBwGXMbJfT3SMzLTJ1x2bUR/0pJ1ueIjxP9Mjjnfolzwxy
zAwlktVw8TZ/p1JCQ7+6oek9v6v+eq5WyCI703pMOvlCBAtRBu8wLQ9sMRNSsrw8XMO8SX6Po/5Q
5YtwVws6v7j6RNqU1HvH6ZTSZVGu7j56kJwhXpkk5pul4gEc6RyF+NmJV5nc6gz5QUMdvEigIPxc
ECtw0b8E3a3Ey62sqln58GMaRTcyX2ghap6/1p2lCOzQdo+8sTQiieU1jjL+/I3e6ALYnUVVRxEy
IxVzXBAq+zQbQVvQDm01DPpVTaa/ThpUexsA2/xSKpbQ/N6CVjP4/zcmiGATrUiAHZDz++59ehm9
RTzhHWsn6KCZYfwtl8rAI79ElzcMcEZNfH10nMXYfADUceNuLVCvxHcyCxK9IhtgFVAs2U/ytpZY
7bXdgpG3uQ+SL4OxWIOUFlj4PSYc545S3SY9iwbHmozbARN8FwJJO74DAEZQMbRlBMLQsNgXOUf1
fy8kYHtJlLFoMCTxVrnlo4DbUZcCQZrHoScUEDWtBPNJEzOiprL12Hh95LNUlCOeDRTlSIVkW8FR
1+s7OR9aeqoGKU94Xvc5rlVZA06MiGPvwe21HTWW3QVxASIAWIzQlMZTuOhRZCyINyW3qcm4GOna
ye363LJayilFJRe38UVHuyCjP5ol4czmLGFtUYMBnFk6ab1IAdeJOl4wbbWKIPuhifFbGTK9YRQa
HBz9bo/3T7ny6u4dQZ3Kxb55JlMnxI5MZfUVTL9qvH+smC9rYm4jNF5ZazYb5jOdlj1Mw0DRVHjG
od5H6rOts7c3U+nkUPhDrVqmVcymoRUA6a+DNyLdrTFVKEVkIBwgqC5yA9LZuvQD8vX1bwG2FKtF
MiktIolnfF12KyFt/1sq2HV8uL4wiMHQBdOjypPsdcUv4q+df/MNiv+gcLMw4zEPSX3n5qkdL3iU
BUZTlzDv+tvjzNUvPWYGzm9avmRCtiEE0mYkWByyGNJQm301M/FVN2eMQbeWCVeKiV2/vtUx4qU4
4KqrFUrnm8EF5mzCaI55ITGeskKOeSCETz6NTAkQ564LGcqF3tA2KFfZdVnFjhnaNsWTlJzLZC7s
Cnhi2NeFNuTJ4UDwL/lWFudJWa6EPEuilfqA8bE3A2e5PUG0TBb/PSM25hncIWBK521s8VmrDvkt
SuoJugxLChORwVhvTaLJQXx4hEDtC7Pvtms48OfWhezFxx086ZI4q62PmjTS012q6zuTUsRUANmV
sKYAYi3VxyaId0zw+HS3npsnbU6oB8Vi22Oa/9X12lOaHIFhauoRiP4VyI/c78KULRYDMfZIK+wW
4eY8DYrtSHW9zXCsTVwuL2QrRJA+VraPpTEHWmdqKGQZBYb9C76i4BsfRl/ZtALkZ8FD6TlzAIvD
XJT9vZ+5lTbSoNVv1J4KcjU3mDRCcZRQIa/X5092DHWGeyG5EceUf9evwiJUi50eBv7bao/sJexf
GRQL+UcQWbN09iyKfz32QgPKj9VrtjbbfRLYalDEJpPBG9bmeBWSMJiyu7A36e9mfDcT/ODWpoET
sBoIAoBTAB63OGy6grpQK11gKZCCPMZV8KONkHjgHsK6kF5Z/wTyuK3AGEzmxHmsTTrbRk7lHIly
4yxrNFG43xMgLxJ59eojCKXbR36DUxpETgPH+MX74lBi/1HFrf189m8jojFFBeMy2YvnhIIxZI74
+LM7favepzmVe7LZQRZ0kavJ3emByZF/GUG3Bwo/J/MpeK0rxzFjKJn+OkEkV6ZcQZdJM0uBURPD
NRM2DQ6oI9cg5CiE7oPgB1ZPFOoWPB098OeG7DoMfmWfPakOP+TgzKuml1iC6e7SrHnSx4k2V+UZ
E9GWgU32jeABTurlFubIxhC66pw6O2CrfMq69rd7b4z7FKSIbcCNd62zosAUcLPqvpv8JU3xMqIX
KTKPWeqklB+HA/gKb8PnjOZfSKNGFGrfcLWbm54NlU6ePc3WRlJ4dVUBaJgpmW3FhkgTxw1xd+Ip
PVQxBrVTFqonbkD0a/gSYOe6jXIQ2JWv+/iC/meDHHNv+lkB4YJfwfhbIQM+rEzWfU1Vjusakmff
UxYYu81XxQ3MseiBCW9Ei2t/OhAydIpFWpbdssXBAyiJmSK9qHbfKeRvFgfEvpqZRTk0jCOl0/hO
92HH2dxZRBWiW08YRTdlKcPlQBb3o75BE4ALZnEps9Ja43FAygjr8doQaHvBSBbnRAf3mUXzz1YA
QSsapqYaqN5+TMVk7anmMd7dcll5QxaB7my+k7K1msZcsOMtQql8k+cymhiDzI4KEWbIq18q0LEz
KA0b5atHcEWgCGj41W4BUrJr62Q5BRNn2FCYPksYT+bwGXXSstCMAL9WZb0/bU7tG0y+nRGxPwbc
VfToi4UmwThi3IlM/CHcYHPFxhQl/NHjDmr+lMTinUDEEBY05xfJN2/0LymYTKNkQp+caHomX4+R
XWWUoFf9UztG4CO5xgLsRMZ337LOarlFFBX3yUWwzYhXY++LLhUQaL+SZ5ELpymhL+6XIuH5XF7/
/Z1PoNofoO14DGcXYaMrvi0vN5lh9nTmyws5YhnleZS4sr8KCYPXT1M0kjEPcuZNoWZ4hgAKZAIj
9Mb7iCZhcMJK5ld/oO2F0barduGyFougUunYCiCgZ7VGDjcFB610AV9kieSef3DFFfT6nYXq+Gnf
z/m2XREKzlD/41K63d/VpUx9GsvYT2Dw9mNXMkOnJSqCCRIlbqIK+VGiQ53CcG5zuClk4/v0HJEs
coiwMEq86Wb7CQ+O9QvsE21EipzCfDS8bkTE6iaw84cDJxTcd5XhrZYB7vo9NlJPBeP/pH1goup+
fWUsIkH6nN5KiVSyHmAjuepUkUgmdQl0HEFSG3IEJXD9yaH14ZuJ1gzsJg7Yphuk10+T7lxCPGEj
E+0HIv9VZyRY8UTqFCNr13DenVVE/aNRFagxtScmlPjmtmgHSbCD2iBoly/7HxunSpr3jH4BHzW9
DTkC8imZ8ybHnLJC46oqmjE9zjneAEr0qlLXV2nPuCQ0+eeX4/m0VCee5I9uNeQFULL0oImXgMIk
+Vm2myXYywl8Vb+PDuUCslxqC5sW2STsj4LutEFY9jTPSM5oAi27+CLtWSBh5syDuqVi9tqN6j1c
8JvXGuZrSLSFxGN8yi9GFDs1rNINpCvJSSQ1SxppTnkQgXjBJdBjMqb7mi/TBCAk1geV6PdCLrlW
8GdFxuF8FwBpcPVOBchqV7kIRgxvTtgcP98ml7bhE7DDCbme6X0F+ZSCbqdjTbJPqdNyHBceaK79
4vZfCHX6UY7+n+gCu0DcKWqX/gOwZa0qVlXCVGQWj1XPh3/DQjtIDVQ5sfrRu5o0N9E8R65DqxtR
yqJmf6iwNbuoJRkYc3nGy81ZTic4lVIsSBeHN1dRFa8eT5uyQ2DPwKtN4dOCgKGjvEvPaa31IBRH
WWdeC6Tt3X/qpTQQn1cezb5ydQXxz/RFV5BaziqACbTI8NgSWtqTHJGnm97Dx+ffvPnp4P18vtp4
+eTIcpRPin/g9vc1z6TpzAZqpeBfq+MIQZ+mN/YtJlPhfdO4havOsFZ9WK1MqWYNmrfmyCW3xh4G
UByX9EqUfB3rH1o+V6nRosU3Ub6AxBFYebQgf5iJnt/2J1cH2EqOyOWxLVYUOSJEEhrmK7aEEb7y
xLGOfQyLZsWsvqoRW20KwCdC9TAvEMk53XeVSEqXpMxn6m7DZfUty0pZW7MC3LE59GihAVSiwdOn
1PSy/mvoA9R+qZAXueYNx7zxe7I3yQ8tLyNVQ0B8FjgFu4A20/lIkdTvlJbBbKR0LtUjtRtnj9hA
+co1yqZXxWD4e7DnpeBHJWbaFJSFDQXt8xbMs1LOj8zreerIq0l89ZGTAb/iljvGBSD/ciH6WYo9
iCBNEcLjmQGH7VmiWB0rSgW2q9/Gp9h/wvDTpsCGulVAAmsH+alGKxe/O/hygBPowIama+vc34fc
vMGGfRIDpwLGbT5fzdhvpGiQ74ZQhfqooP7XlFFs7vl1DczULp3VV/E+BxqiXI7XYqFyvjrVqVEg
VjuJGAPPQuhbrdGyKzCJ1AtunDjZ/orzlwwN0CtPXnW0Ff/KFJjT6XSUfQ5DN8cDIVz/DhIAMyYh
hQKYjqzs3OFdaG5UZgUeJrMubhqhP218NHOI2qgmrfdIKhyg+i/WPX5aHnvT1vhrZPAYueutI8eH
fUaEtFKmw1wdW6vZdmYb8KCmTWI2l0r8YdG+fUvlxsrMiRV4ZCVDFRT1TOu5IWtLdRNZeHXHWvNz
Rxt67NMt5sTRJvlSstoSLyFJMARBVpIpEMv435LrwFK9wHQttnftyNo5HYPlLzvyhFjQjlad64e+
7xSd5B291HDIWA7T0spC4Fz5/Dpfaz7MvEi0KLfHvvq2Jz0K3tu2V6XldpOXLGpi2UDmmFs53iYB
+aUk60Cije/qBr8HWR+5CjNecVEDDJK3B9HOgQRgs/gw7ahBtVv5nAiA1evNFKGHK8oneLrqqW6i
Bb2Z30E4gqDn6kKHEzBlEmHUYik40eB+YtcNZJXsDl5GUqOvXclhAZEAWGC0vJLony24STqtUIig
pOOLtoPvwnES4xWbF0MQPjsUIXVrb2MOPM9ivsKib+6uCZlLRPTqq6BJ+97CB+6FhbI3gLzQdpQc
nusZtWRWd0JwtzzplLihwXWy7+/J/JqEMdctlfE2HYHrT8HiA3MUXR7N1ly9xSrnCaOT3/18P7Mk
ucKFS+Y8TVADFnvk/WTOQfT+hBXEXetc/rFuOlicGnm1e5+0mrbEQaSriBKRBj+cr3rnFSltoice
NGLGQJz+qLUYpFj2tqclTqR7aWtqGHJL82eYNZNwVkW2b11zXeFMhjRoeBl5fEX/5MJWyigpWRJd
wJkbA32ULIoGnXGW8muP5Osp6jCEcf98v3K5uQmXO/xsIC/oCVs6+H4bgrc3WCtsturkkNG57Nqg
cvLS3BM+PFjhWlEOCaM6w9KIlVKheAfvvsVW6uM7742TgIuDg67ijt+wGRsrjy4R8OKAUXk6d0fR
1NkxI+ZNuXbv2gYlur3CdLdqJ4N+rwk9V2pU8+jg4WfnR960mF789i0+R7VrxQbtkPtb+7kt69Kc
xdIMrfnLKSCOAMgHeml79gojSb9w/b276sOCjtnleqozqko0L9IL0swP1Pqt66wXyvch8ZFZ5Y4o
Z+DkIqaHWFM6PuP96EhBr2jxrROkXkfkkqGjjPehVt4crn3IPcB/RUWtT3mGyEcil2VfpnZCeQqy
bb32jMpNuXJa2xtNg5brbLkvX5Ttcf5ieX2FRquGRn9I4YmnzmN9wuhUHQ0IRKrMxhsCmqPc6VKM
ta8PWj50J1qvoPydGjt1cP1Z1W6V8Ndn+QtHwozgkvjA5eIykKD6rxFLPUGLRKyfW1/UgWccUVk4
ioIcYVWBlwNdozTGn2PfRx5pdfdBJB+MtrCCsUJd1mElQfg8g1UqaAECZD6Z/232LLoXs5idnnUi
4A39FeqRzgSfrpVnz1v5Rh2JoOVvrHqzStiEEGVjPUSOJ0pC4gAzRjReps8uDygH2ro018iKpJZW
KngcXQ3yqrolKm6q6/Ny9Rm7yqLMsznQlfyN2oq4xrcKa6CsuuoWyNbp6UJGxhLQValmUoctAeg2
/VF+26zwG9uhMh8+0exDgHxhtO2Lk3b9QulkdM4ubJQ7FztakfjeYnSKyA69KSjmsH9x0M677Y20
1xcHEaOnnfKfqG1Xsv0uUN27ouT2yMIfXvGrRshSAcYMQ9x2xsiOEvhC2N6ibTDkpeb7kEDEK6sL
CZAlkrWw3D8lDvAyjI/n84wxQDz2rxEsqVPxbNhTYqesEIFPEw6Q4ASYjvjy11+v7iVoeg2UppgH
SFjNUXMcUcTFQwzMDJKF2sLxJm4PTeL2y627f+7UOUFkdsx4oYKdWnhEKvL+1phzfXF0C7uptUG7
mHa2hJq2b24Yx2HI6l9Yv7C5InB+Nytfrdf6KE9QN8J5aCXcN1ZNItYQAlly2AZl6LPN/QU71/Mh
PRULb9i2cBhKTmLeE4/7KYbfRkhRG0V8NOyiE/z2WnLjqxpdpOR5kyJfRMWdY853b5LoBq+slWuH
JcnPvllGMYVi98BO+ZjIQJUvBHlH46n+MGe2UNNObwgpG1KzKV1Xy8WnK4cDmlLgIv4iEM2mkSzq
56GcMnmmP6wi2kFVoDcrrFpk4PBZND8TUzMHdvu4nDOASN7KYQ1VBotCTyCFmX5Gk7qR922ASxmQ
zxFgexUJDjjxJ1Lh0ve2O74OATDEXczvnwHJElEeEBdrAbhJH4Zwpvt78yU5NRL/cCJkl2cQgfli
zvoViPGBtBc7SIwg9tyvzHwK5YW/v3sS4oU6bE8fvnEUNezTFzV+NzqqnTym3s4ThKiaIU2/yuyf
io6VkFfeL7bXVbfy2N7VpGDRWr0l+gphKc+rQtNLgIFg5F7CNMQknVEOx35JL8Lx5uM80Gj07vM+
xsIc/PhEDsD0SHEDyysNWJropy4i5D52xGIOcm0+DT8kX5kejEbeGLmQr6PgXmPPb6oiwZu/mFek
Cz62TiL3b2pX9evQhaskZm+x3dZfqVF4n1uiL9nLduT4h72PHNBh+SXrIcfBmcvEFPbJ7oCoAttO
i4GgZMllb6hBHxrIWWk3XRTRCm4bMhDyD0mvCf3bZ8PxAgGz3BNwMIkSjp3dRHue/Bk5oZatJFiu
ja66DO3haiIfd0SGCHwOFdJ9LHS9eFGoKFK3PzYeNbngDo8vXdsQJJTNN0jvn3RASKVlk/W3ZKKU
xvHhtSGMVh3fLf5GWPfyDE1NgNYqG7pcMmLcKkgp6d0UkgB1mWIte+a52y1Uibr830Yp86Tlu/Ys
AEuEUCIgw/SUppj490p4yU3yZY8tH9Vln1oCDAYMBtRhpJLDHiGx1U1UQXUy+Tb8nI2sDTqV/BZA
ysj7YpQUbC8wTA61gyOzX03/QrryHKb4lqZthee9MMFFan17ppH3WtA7owvS2EAD+UVuRKCwHq04
rY2uV7wYXVc9tD9tCpuWh3LttAGYhRxSgfpXb0bj/dvGPluYFKjJAq+b9nYFTSIvF+uA2fE91P92
xpXeIQTNHMkAqLHW1M+uMZ8lswiTv9qswdH1Qx23tTMalyt2GkJ0j/d1f23AXz90RoNp6sEHqEdy
RuxyBq2CG3P1qY9jO4/fXRD3yTDIbmw8Y3aPtx3MyjtfOdQDfI/Lx9zYt36gnippkoNNMaYzB/8r
O8IN3k990nrzbN7gpr2v1swUlF6p3nT72FRswT1T3btpZQBuIOoFYCTtKzD8L5LPzWKRWDxzfOls
T+DRPsELyp9FI9XOMr8JS9VaWsp/rTFvPvDVCyk2to0ZfhUA9gZWFuV6zdf922Te00MsU6PcW94Y
CEX9P6QGp/T3ZuVaC3ev76SqtMnW5jalTaTDQdnIA6h+isji9KOpa5B3QMtUPywKzymX7nmmsdoE
qwFpugusRo7RCbaZp4qJQRERlueGtDJGzTosnAitRZ2b2o/wHO1SHavcuAmLzXUON895YeQlamd9
mQGXdDLpmm2MLeHobTP94jyQNJWqCMhwd9JvN6f4+SwDJ6iuPezEdVvsGT/P5qXXT+f+Ac0RADnx
OeCNQRppESan7JN5y/QNYDYERA3tc5+AJEOBaO7kbq8/G98tVexSiuWA5LmCGSUjYB1jhGHZ+9hx
qWAHNxa6a0OHk/6DGkk4RJtSH7TZDeDMAcGpXqLe6MSrcIpjOKtSnz37Hw79VG3+bLVUuHAwEfrf
D4GvYm2VjyBor/8qDzJ6DbstIEgKyRsaFy0ZMi2NxMGWqyXnA15uuucWj/sktk7PAtGKAzbkywiV
LKYyj8x9Qdlv0xhOHNq0IoSAf6ijpAK+xpDCp8aqoJDoPtuhZMTKeNd78HGz40M6q7wpJYug7nBz
f/PIcqguL7fk/bh5K1NfV/lka7d9OA0yxiqCvFURKdyU/6Ge5LhO4N6f5nTAfbtiwfyic1sd9x4E
CSXY+OxOmErBf8ZruvKt7pBVm+veU9hjilyHlNHxmO82f9IjVPEPHncH9rEdkc4QPT3VQTgX+jqz
qUlTaPHvPaOMP1aSnsF0peNlb+M0jNTp731I7q6Mp5xnN8WuODXoVirFzNZzO5b6SEIahHXHDSHC
LApiBr5FXovV7LeFfr/S7XdJFUnnZUC8tjNCEsZnbgeQ9Ko/NO5fT4PoV+z/lSRi/Dxq9RLEBqul
k3Q5SLOC2jZLRVhgx+xzAJ4G5ooK2cGQ9aaswSby5SUQ4z6gsHZj0ssBrb8fHdWNDsIUGYeK/2xf
20y/cms3EcRAyR1IpBBqKfTpoWJhVDw7ApVqXK3RrnCtvg/eAoEqadDS5zJGqVzp7wVyQqRgQQGl
wWG72ZocdYPJKuFfwItTEhxzK783zrgjs7LwZAVoySxRe5Wzkryb70ay2sqmGuAAEHFLeL9w+W32
644jlN/ZAypzhqpqKqsDRM/RRQcIIkgH2heofgoM4EjEh510+Bt1F0d2G79QTUr08IZQo5yTo87o
koq5p0HDfNsjH88zdA/J5hnsE0ALuIcu9jS/nOkSDfq2aahBF55IfnoJC0zgwhBCR/IrEdBWCuv/
/RXqRfVP3SabxpBnDeoONZ8hzgU/H8dUoVHyKTMqVGOeue9pZnH+X1lx4y6LAeC7yGaqlVL1871a
0JGAEExlsqTxHs/YC2/uZQQvecem3TA4DD/fbz1UgsIeYmiRoVjfU7CJCMFJY6N22EbD6M7+yaZk
0FHtIiKbu8htxddCHQ4wiSd8koPeWOZirAs4mqGTqdExoEsew6EIodPAHo7B1O1DHY8lmFw/Boqr
reCUHi4sNLE/Mae3kSXicjVZx2BH/HlhZT1IbOmFivrn0VF3jNiKEiF1CDuEtnGa9fikI4gpVLO5
5gqJgP72J5f9R5Tg5wnwyBvI4wBLmIFVHUDTza467mXzoGnNsFrXCvTmFpEqIY//pZ16hsgaoJR0
1YmMCvlh2m5s9ViMfkq96oEGnwtgslzZXwq1qR0MqPZKci1Anr4VxElVFCC3z7Oohin0AfHLcenK
IOkBAB152/POVFDbnjiJ/X6VJUgArGGLXDPJ6Qb2ZBIzkcgaLRp0vObzcO+K9h+uXLjPObsxC0MN
NemSqC1OfskurbEsAT0Sc/6IsdI4TZG41BR3vXg0c+FhEcIdt0ggTenmUI1TepZg6G5zmNtM+NwC
nzitNxPKd3nBswBo486vs7a4XekKKbEKd7T9/5J0PVzVQZdZieNqAu8YCQ0Ql+wjt6E3qsvIWDRQ
l+6Cg9gOVsDynnkUgbTDW5zSGAcqz0yKVagdZ3PsMlk4sQ6Vq6HnWdtOVceplFiZ9o5oYCeonm1a
QurVwYiweDx0N2G28U3YFanJ0BCTDmh8jsqBAK4Bs/4+TlBsYp1qm3+aYQ3nYNHJg+eaDsGlYzRl
nbmBNSDxOzQ/cBB3Gwumk7o+kj9sjpUbQzmpM8BPuHHNi1wozVu7E/lfAe7ZibYgnkTvzGcpkL6w
dHgrXPVuJo7N+43VWGHVWesZFTXWX8EQqc4v0XpljLdykztaH3PeEn89SR///8FhEUsFnKD98sL7
rVnSh8rK1QwIwTRdlR3r9OC9Q/muv1hL2jqDScBPg6tsnQLACFZabTtbGFzh/KLUmKVJg64k5shc
FIVmaDHXbBNt7sSUKx4yTY3AdoUArclhAGq/8ITnxvkK7nw0uhDhNO2sS2uNHdp5HV2Urr8IzWx7
CRaAcTUNP34WY81nT+geYav8RLUvVmwDLPBIjtYArugUXr63YIYu25d0Z6Bzz+RhnQmLjbqqaUGG
7OF4LcKp6HrCNkGpy9IhefLMYRnI8o8Mg0vXkiWoSsygXO/Rk9SovHC9tlLCql9PHKA0wkESNiiL
+IeMGsQ4doSiEeeCMEG9yHgxQwEF6e/6zxW75cKTmREUzF+7A0lThnNAksPTTRie7SqqIiLSrjcU
YB/iCt0lbjczkxJDSMLtQJBAtxCqFAdQejpTJ/b3My8q0GIrz7vlOETsPkCK6MgEOHt26NHy1w00
YTPMtIAXOx2uUS612D0Q04NdKMjc2+/kcKofp7vyjWgVgfQYIHR1f5QGUL7Jyvo5HiyQwKzl1Cbt
l95HepSMkcxgjT3VWCUnb39AFREE1qNYzdJR97dQw6fLlYPdLGJFImMFQcXJSxlvHW6yVPxQMtS2
VjJSZjpenPdfsNQC1HafNasnFtLpC9Tkvsd/sYC/tQfU1W+Rt+b3XuX25mxfr0U04cri+sOjuUb9
SkKjlpSJthrDWxj+6AmR4e6X7ORpNEz9bxyzDmlCl0H46Wfti0wEx2j82WHa6nzvBknN6U/1sBCm
UIFcYB6EIC8ajPT+sx85O/nEZs9oUppY6xL1bk4tPevaHLu8FmfaoCnjTYEVBFCPj77vEyWF6aRi
1rz6+FEnn/wfi+peVTWwj5ExesnrrjNLCPB7vXmWhHz5WWpduy1wOWzz31D/zBzTQvg71J5t8A1h
nBUNM+MOoAs+mVTPdt3aummk+VzznENRiHxSadRf2lFyPqmDdMTJ6W0JgH18l4omm6u0WxNMNB0b
tpCcoDEH1F4Etr7HvK+uETBg0/DZktrewOvfLfvbQ1OxqdrngNfH5km8MBorT0tSHT/SD7Mzsy8n
2KoYTcpCNbbP95m4Fmza5exVLwP9M64Q5ttD6f6OtQKnOL2VwVkd1Ax2ioVr1z6MI4hxRPYNStAJ
uZ/WDCWA64BdwFtq4OeYHrdtIdukvgJ52kqXwd4kREvOE08RJPLXurgZlYRd567I9s3FPUSsQhCX
/4lHw2Do4ZR795rs5wUstimBcwGsy4kBny3wn1Pbum0eb5bqC9CGHdLqsHsHwQR/b8msYr5D/TK9
Rl1z6XJ6epFUuHLiwedYq5tSG3Gp/Jr2NJW2M8ggjdESUR4ELr+fRqZb14tFkd01mzM+AQ3ZyO6Z
1OH2tfcSHmFJ/FYA+xqXrsEstHJRujymfevyZp28R5p34FYsu78l2n7qhv8qJeof+/G0thtD+Mqa
k2AhPg0OBMohZSE1X6lZkUoFaLGE4FcmlSM8g6ANCAnuowHnqHrSDBqvfvHg/BVEP1ewQPNCjL2M
SGDgMa9BuNf543tW9/U3v1Pn9JveRYIEa4Nt019A7wJG5GheCiXEm8cEwyAuIX4X2S6sr2VgkCPE
o2NfD+lY1FHzF69PT5HLUnqDs9RuZ2WWRL6zSVsGtTd5pAnmbloneIOXn3T5htZw7JhDbxM69NGC
042q1Pi0Goozq5BUamf/83DNs1FI/IwdO2a4flnRToztyioboKnpPd+P7tGIi5MRk0QrVGul9SyI
xIQam50oq1k2ukIy7onWztrUSfxGZnWL5zXizPJQiFJDKHnAoKBtd/17OSLAUnYgPkCE7K607dtL
J2S82rgyVKwyyXYmeih+nDQ8gg1C8cV4qJavYFeCAeV813+6Q37XuhwhTfDYcL8laaMrKv48sgfO
ve+LVdfZ5PnfMFXnu78c9ndaCO73QgX9UKtz3h2ega93AFuFYiGuugqNfhYtb9QT+ByzhGanBvkI
DJ4Sq2M5n2SavfihQVpDVN3XLEBhCdxkgMyQvCzh23LB8WQK5GJKzz8Bkg1cVcPSXL8MGmmH+yzq
zO9Pk5+byS+gVobfaulTYq+id63NSnAN7UhAMLJ7M66oK9/uOzRVrcX8KaT6VNNtU+ejftf6YTjq
ZqT9+UWMrDyAXDDagJYS5b60yA7wrNtKYYO264zOThul1m4ue2Vqe92VpLgOBk3VfvdUnI5tBPuA
2AbTJjFOzeT92Ws1rim8IdI+d1xfw+KUeJsnMjZf435uXLB5hNLIMY0ddKk4/d/lYRzT+ibE1Os5
/t7Pj7/BsWrNzSxZDb45xfo9Yy+2hS4v4KkRuvWnQ0c8WS8KnfWy0EO7BAO9Q4TrcWEIOS2G7UhY
bnB2ONxfgk0VcS5et5ZpEVphrreVZslvv/5co3Z0DI/36tlEDJRUgRHVG04sJgQIK2XQqUIhSvGv
2C9UGsblCDKogR2oRaJVBYQMXAJzY47jzyoijrLcrVPwOZAa2kiWBKhyQ5vtpZGlqSi0nd3FAM/U
XrbpM9XEgYDOeEIUitaa1DpNVzP9ojfZjkVobpeTt9pXsB1n12EOc5P1Ruy2l+N2e1NCbPAwSoib
29RtPJ9rBlKagg29Tt+5c+AeM5bPY1UZYEeylznfoEiwabmRS39YV+6Vu6XUA6YqyiHEeBpvxyoo
oIPJBnEaoaen5X1s71tJpt+GHpYT0TdJgQb97R942H/gk082aTXfuIuOP98eVkQjVbIsPvsbw2nu
G/v5nk3D+qtTg5WSshZp3+4+p2iRaen2mey9UpCDlAs2FqQg6Fz0hSHrJvJaKVM/dMt5pFYkRg5V
dBHBwgMM2mouXUmFg7p2LrLL4cLh6xIseYa8fHYxNH2K7++6Uo1AT21SNA+hDLu+6yVAwrHoecGK
5HKN7e3FwNq4DQ+64eH02TtRi8z2pcYnU0C5aFrTiRI9fSSu5jOJh5oSUmFPBwB8cjS9Cs8g78U0
xE+nBVzKCat439Hy+BNhjZ+Z9CZL0pDdcjc46GpBvzCVS3ibS0Vv5BvkTdGS9rakNvc9LLh6ofvs
ExTQm7J4gNvS+UgojPYFwTe5yOzMVldx3AH899O41UeWqddnI5YT6DwBudEWpPDxGh5pIRl3J33h
ovOcd2/ZAFFtSMuA5y+DIHjfe8gfas9lvtcEBMyeBpYQvh/+/hLyEJbKopmxuxl4EINuXgLBnr4A
VmAUO+MIC13QcdZuigB9NFOkLxnj0ENlmwDYQN+Wu8J/vsREc9Lvx6Mjy/kRFDry+jVuTinI23zt
lSoXRD2uWviYGUcoFActOb10CwSMFs98HItR40I1YU/PeDNqUx+6GrwjkbI6CSNe7Ddd1ld9ynrg
4brZaQKO8ILzK/Hb+S3v9tJdF4cNv4kt1o20aep4zxWsXe2Ih/c09qtx2PtjHIuBy2TfV6p13ihe
1y6DXZ3VOIEmPDfH5DwvcALl7ls5v8IpVYdG05LIDKBFXMdEM+IDZV62sgo9p1j2jPFI6XOOXrOz
Gi5yqSGVK+0Fgs5J0FD+1PZsMDFlh6tzQ1pZqd+tUJaM3regKKeETRdRpL6EWV2GjWUym2O1Sm4h
Cw4NCvODdH5KtvgvjGJVcE+lTpG1r+rh8haom6IQatKJfC4QuLIu1QQNZU/l6+V8gAOfU3j9XEyC
30gsnDjIpNEio+auys+dWTdDsX/wf9nfZRNnJquU9sRhjazn64BILl1QXyIf4Zz36Wu4h2frhylq
hRoQsJcgvHshn1o5nu0xX5tas3LG7f3GAZK9KW7VpmslOVV5tz2o9LUJz3P1BCLDRER9WXRfwigY
ckdFZdxYdnBUuZEQDSikJLHa49FQB/AJk8W0xP5ojtsbqlX3r9nqz2De265HFWeB4kZI8SoO1jvy
fpGk9bxbOjEm0qWlpQXr7nTNmVcvta+BgskrjRGaoe/Oi0KFTqnx5cCaK7w/4yxfkVXUBMod3Mah
p3L4I+ykSXz1WKtLszmObSHk3Ca5u9obf87jEAxIJvNxIYT7L+K/354n2wLWnvcsbWy1xbRx4qeZ
dQ6Yjqg5FCP9K3jSwSRYLxWnH8dE2m9KXg6gV/pnYy6FIcToGk2msTfO2Q3/vyg9gqcc7mi+T4ay
qUYYjO87oXp1vEPJjKLoIuCxqe97C+xSM8ylybcT1kr3pb6al1PLj6p2n4RPStoFp2Ou/U736Pev
NnWJlmAmazonZVSGW0jo6svjaHA0THR7opscPVJQCM/gbtj8RIsOHhP09PE2CTjfODmLVLL7dllk
kfdrXUaSAYvmnSes7dH9AwkgLjn+MSTmtst6Bx2N8cQbUlQ90s1nYhm7jycVW2U+hJEMoEZQijBm
pZ9KkmP/ZBEpPtVdV7SlCLo/FNY4ZBcbRjsZzMH2tRPTJ3sRLcnzgMi6A+Q9C7h97EWogxdlGkKL
1p9Zr3JQeK2DN7VnA7vfsHZ0+H0T/UbovMJPBakEic7ECzAbYMADGU9fWrKN1SsZVIDXaXgp5AvY
oq4l5FfK+sCu/s+N2e4ISlwrxnO+qDNV3+FjdRNbGvBaP5MTfVKwgOUeP0TPDF50vDV0dZTx3yOp
gKaMKnYFcxkbxN5IXDCNWMrICDwMlTnYB8ZsQOCLPorL9CXQXqhs8cl3Iyc6uJX8n84OhZ18Or77
pyGYIOakmbQZ1S2lg2zoS6o+EnLmILU6dr+cLPsbW3lu0xo4wQdTCOd+Xa8izfyah1XTcGQusAYB
5e9a+9z7dc1xJvrdqWzswaFYnUhbiyb0eWCrkmBHblEMTl/QK627hiafmCMQqhxLr9A8dGtAhbCD
i7WBwJJMMNuEepYOJgxLmaEbDdw+vOeHlLo7ehKva+vz3xL/CJZ9ChVJPrNzpejwXAwd8ifEk4Tw
6WnJw2tWKo0ye7BH5sjZQXXpmyZXgXcul5zG3nfC/d1vXB84zJI2ly657xnoaHrtiOlLFeNaKLVF
WRa4U9ePUtohNT6c7VM5J6EFOV41jW/Xx5giDpkLkVOnd1XFyPeyArxZ5jLy+GyLZqkClflfFPf5
Of+dklpwOLlhaX+D16ZHP/j/7VyKq8I467rwds3FvSw3sqqTESXp3Bk9XNa3HgCwwUsomftG0Ogu
f+BTHkgp8zLoWvXhdimEGWkdX6dZO1W48zg1yuGjPu+IMLmwU1h2JchbFvhJkboDw5zH1nM0sgDF
jP2kOOq7Wbw3CG8p7P62SCYvEADGHmfaRW0Bd03RhkcFZT1XvZDHjqUjCjPkzRLbP34Dnbmy26M0
MOZ5a7apiNFCjjP1DfbmsOWKufkDyBTcJPOl8AKM8GjxS21zUDYpgWBBwQXspsg80Rx1C2BYp/1x
ThxTfi2kOLPxoujD8ZZk4gmvWquLKBwcnaXE4dJWhsNt7sEqCWWbDuqCIH998RBMgINea6rpXkY0
BV5AA8ayEY5k6SV5xZL3TTO46hqrz+1Ti/Y3OsSOCAD8c7h5WYYnsBj2c/KkoGWpBnZp88EVjMVw
gUQZxdj06R9jRXe5+SDXxY8GrDYtcvL9Sw+jwadK7hJuso+UCt/VqY3iKs3v/CvgtdIjkvx4PoLM
XdvRbPb1/3YVb47tf0RYS7sTj24J0sriIWCg+ymVHY4t2y7IdC37VradN5VItmz1LpMKHE9RlfoO
rB0Np3gBgWp/63C68lMO1EJKIFs2odAmNydclTh0U+GmD/AXP9LAGK821SXCwV0aAPmODtYELfUa
xODK5AE+Tn2VyCZ5901tjT4GlaQ3u7pfXPhhQZapGldUGzN5XNXglgaM8Bxhk8yn2O7Hn7bCrf6z
PcBhFzqS8WFGfHacI1/oaHL7onIWzLAUJrBuBDBLuiVjeK2mpqwRHwSgqKBfU0cgzx0uqwxaqSe7
ylPdTlhM2c7XU58weRxbqpvABGeClRMnx0Mtlf2IppxRoMapjWsK8n+nAzrB89YEmJJV2C8J+rjC
2hU8AOVc5mscGBItKaHLKy5e5lc9Pmy8nelJmmji6qwQVtALzJ+hFXUnWCqAP3GIrLbHVkCEx7xF
NXhxA0PyQ6j0kyZi7TUBSs02Jp40hGdyHxrZX2DkVatEV8b1ICXh4+a+J2iqsIizSev8cvZtXRjb
5f60q+hq95DFuNcEwZPqVbfQQSr+/x4jXAIU7IyCTo9ZTzyNgXXWb1DLyyAINFV8f9dQKE7Md1VV
JAskgaX8psO51ujAsqmSfDVt8Svdi1meGAjaMWCSMIz0g9kDFYa9R7Wfa2HtmLS8YsZB1nbWgvbD
mcnte7VO6SxoK/ZEY+GE4/vRUCDSX9KLZT3Mp2tuMpV+p9gJYbhBmIvLLILGRA2bd+h5E+DnqMqQ
XXpkBfqwARPE/LWIAauTp9KuV7LLoDke8NpkruJx6POve1EpUb4LN6Y/YMIqsy+cBr8JybgbUUj2
vxcoMsYb//dHYFP1DGRHX4P4MPEzuel3laODdYwznfRpR3vkVtns2TI3U/QefgojohRzJj/UXs+g
7SzcfyEHGvddj0SzP5/Avs2kltVHPAK2YrLAdDdhiEKerKnWBnmwHGDLEoq/Igfl7yvBz0vlVgUh
UfaCW0Z7RijdwYZDKAOsClSdev8BS47AsTOOUelGA4tMVQYBRn3bEUxdCHHmwx5zAg6l8YUOjgCs
pQ61G8ajrbuBfIwDwvvidvcirdvPih6K4+ISd4LHf5J9S8IcMAPPwbdvyoteVEgJUvZeBCkuq/rA
JQSiPqBqLRV8Fny3kF5HaK/KVi6LMqVsfIdj+7fcwTrtlBf9vQ614K1NgVcAaUy/ExhjiWw1o6T7
vpymDwVCC+jFjG11aPs1wJl4l1ya5f6hHsLFL88rkFw1DqbwBF2LYBjLjIMMRVR6N8snqk459+w1
5b063UPNtqwYstJyAlRUq+KWuXPSEcAET5TZV3RaBVdodhnz9IjInOeacSrpD0Feu0Wk1wtqTbvw
0JhID5W3rfAtNPbzLpgBqciGb77qYB1P0CnDkTkGtioFV61ZTACRjzRt0pqZ6HYk7PWD2b+jAhaq
1jClNSzAOL5/bh1WRc/mGarKWTxLNWxOJu/MW3zBbqH+0nwIt0ZViKIujUgshL1/Uc4gh4r1Bqu9
21Q1jBhfKJwoxW5Ha2Oj66Sqf23O40NL6czp0zsJJSuEu9FlkZyi7PB8Z1WeyE8pkUaMMAQfGa8N
5y0hsb8UsGURpCKHaksgutq9yzar8YMJ/jjrHk9hbgAPdvDcnEsF9x980Ls9qmOvuabqv3srQNy7
v5pJPX3Vi5/FJRyxunzqGiFWOAQiUD9zRETXKfmY8VYcJ6eyz8EZLLqDTJbAKFEuvlpyfHlI11T0
NG74opuJNpCT6KIXk4/iw1ENKmpOnqibKBsEnTCYy3O/1uaGOtmXYGEhfGirdpUa301RUfka6sCA
NcMFbjTXeXcOyr/QQQAwlYb4uM5t7I3y2VY1OoVIeVDrPQsLg3CJXj3gaewmp3gNADprEYWReCzg
6qt8coogTsxveY/YSXTKwjFczYdGYbjSF7Ktl8Xr066hrn9tDXzMret6evL6E0AEVFlDN38JltNO
oRImzdIpxk7bgq3kd4h3sqy4O/fByY3qD6VmJCHuzNOsvAPdURCGXgrsY6zAYyMBSqMcw28KoWbe
X8Fkz65jIKvEXXKT9kDbTDciUqstt/aTV++x6yQMUNVTEXBwawQkr+QtfPJxvFlNov6FA4TTJS3b
PiPR+eUPpASR5RlCtdgM8qFdczDImMI6iBSrO01DHZnPwC2k/jHVXwjUKlw0LuuEHOHSTZ8PBVC9
iM+32tV3jPsyU16KCKEhVPu+cnyKutB+SwuCz0mRYzd9vOwPXM7pLGYTZ8mT8hMmJgK2paVy+mLd
ufFJbX6soKFyqpfI0xyXR0sLEMC9X77iq/rZlqAKTPCUsB3XCbQ4A8ZyxmPa+q+5a0zJc53QM7Z1
xLlhSsSKnK7SP2C3oP3rp8b6DEe2tcDIshYG109vyB9CQfM7HhjLxJyuJYkmIT1s2RM9uOBNbBlt
w9eZpqsn0N5zvX+Y/42ZLd2pkaa+16Iieu894x/1R9s963VvRJoHwbbx4KtskRvF5vPvvweQ9fX9
otn0yoQXmWdHDqpEm0t256gcVnE/Da5fGjbc7MZlsM0w47DRzh22uXRJk5p49itPiwp/hC7GxfFH
mQhctOzNtICN4vmwclnPRFyzEYV3FvwC5MGSqDDfXkXhg8Rq4vFzfjDPGl2GVazofkk/v3BljIeU
s8ti7+ah1VrOhV5c5uvP4MJKm15qt76odrqDo6vUZ/FOteBX/prdn8hbqsaigBRmfSbd3whoShI6
m9apGSUjZGkBvuJ/tOn+bfc8ySm5GKkwO3aoMgn4z5LEXjWUyw14OnEs235QykxYdEyBYULZfzUN
kMwYkSNuxuFhgEqJQnj0lhNSz7SdBZkk4IfFQGUfAI0hyDTOpIsKkTL1ysECBgW6pVoHyOXlCAmJ
vSUIGQi6RUxmAcc3ZaZdonBavPIxOGyctvEMZ+QbG878Oz1ODQ0N9OX1nGVp2QygSekSBppGgd3g
KtkpsJz6F/auyAoMEgiTUumjoPGVicX8T8zw+G22Rt3GKlr5gdAZ09aLwVbtMk9F3y0wlDpvpkW7
rrIM/WabIlbzKhzLkleKhO4TxaDmibk+BMEFElyUdpJI+zdJKnx5aeRdHSh6XheClLPTlwbqx7kT
NBAF45TOmSq1bgBCwGJyUwFY74ywvsB+ZoW5pPLPQ6rVoS4aB+2vFLHMetsS963RzcJXN09HgnEn
3i2mN8mQzF6B4yUiSSysvEVAm1ARAm/PcNXG0LPpgBczPIDFR3B8BGndwOpU5eVGa1qLVccy1qsf
Awbu+YbneCf8q8apo8x77J7On6AN92bNjurKHJYpyATuk44lqWwVTRiMFR9uMHxk6uY6wIIwJBfh
U0rI0A0A0zQPynMSmzCgNvVdJIODnlW1W4vaB677RKCIrYma/fCCHPvJDas03QIR9oDuTqaBORqQ
OHXUN4EeAaKUjGbjZdt8zf9qc1KMtK6iZ/niR/DCQH2L6ZLGqPLI0xR6V0Bhg5/yUBhbTghosT+X
jC6D/vg4ncBpmCurnHszaeC95Xhz8A4SbZd8+4YntAhbjlPgSp/sP0Z/Xm2rgGAO2xX/AnwkOhfP
4N/daQctFI9Fio4KlkzX2WcM2U/VwL9AVRup8Qu1C6A9k/8nn/c4BvwSuQ8wwGXaYnpFvCEnE24d
h6IVLLsDs6Y+W3nuHpRbkmyZLBGyZRVLRaghXHTgN8lCtRwqQ3K0X6e19IiF911I+/m6HkLVYaRG
RaV3E+hBjBrnIIMp/Y7xAO4TBPC5aUXKyXHmTu952lae/DALBr7P+Dh5zU8vem/eHetEFcN2S9iF
KwDEzVLMH7PN5cf2+iDCxWfBLrPsG2MgmtodTDsKqw3sasdsu6bjy00kL6sy+I4PPDVnzJbI8QuI
Y3XZs5nWblgOukKxnETRY024ekXnTf40C/4IcpOW8IY0kc5ce3z4l/UyCkCECpOUG9OlRgV+shIs
xIlQ/XpYI0a4oHj4y9QTssjdlolmhtERx/D0TJhn3acQJVqNPzv89VPQzSgsWaDDWb/Kf6WY0pjd
TLQkapR642WtLSg+gsUWbxZ/ouNILZo7/fcWSruwtO2+QjjBQlW7DqtNWCfx8AWaVlZY5BBlDFKs
eT8UUSegEfv8sTGJ1m/+e7ffUJ4c8xH5rP2RysKnz7POVJKD5G0vbL4NRkoDGBaGfIHufvRYd/4S
bISNqX1hoRb+7LKQg5Elut7RsTm/JjCMvznuJnOe1HZ9lL+P4kKVhTBEK1jHTf7oa/EyRXpfHX50
N1ePhNFL5wm61HbBEm0xNeHTlEoc0uFKhOW79G/1N5sQTPxeBULDKxeZxfbsN8alAU/Cl8ET36yk
WeCiiV9st7WuEX5+NKUjbV1Jh1xyLrNsbo5fTtCZT8EPjtzRFS9NNAOBsioMTVZYnQDjtWpKGbby
feEM1Dz0/Eg8Xm3GqKjkJn2MJKijdjANchoBDsTLRLiEP9XMZNj9LVtMF4unbPczG7iqXNpyd8gg
PvFqFaeKk3DVgVGjW6TPDlYx2H58Ob6Rl36xsB/0IPH8P/hWtciZ26qLLt6i03i+q/NiwiuseQ69
Uyuox/aGDBf8sm9tEdKs8eDDgcQwewKGfQVHikPaTuce7NZoqCO34QLJHa9f/ol8Og4z5HVzFxdo
unTrRh8SKDL/yfTk8zmN8JT7UHr9WxwEp6rA6GNlFjjwl1xtI+j8PiHkDxUtebhuxGATJc3mC4uI
MUYv1yb2SJVAbkprvK182EyHxKuGvZ5eTbydkR/MPiN9vT5d59lmI0bZOYN5X+P0bx6Uq0HHnbX0
Swqmvb0Dq22NQIzVX3CultDCBFyTM/tryGambKmL1KShwEDE/N+x1wTNuTpd0ZE4BV01Nf208gsZ
L23y8OLRqmcMJomT1O0wDFjwM21Y257UxJAB0RQZqU9vOkAoq5ztLbguKMxLkN5C8cHjSY2bzaw6
tYMkfR4xX9IJbMqtf/ZnULdpR81N4AWJwBNnW9XZZSk/slqZ2pB+wodemkoeUKcxlQpOiO95RZdy
Y+upSiLTGqGCpbHcv1NMjehe8WUfzc9nfyv6juxPoe0xa+J73cNHDnWelGditJowrlL+nrcIq70f
fy0TNjH0LZkbw7oiOXC9WTX8y1Y1yadRBIkbVliPG4+TzIl6CxdYfle+ACFaSPN7mi4VqcoLWgtY
SUvuzfh9MG7I7aAM/Nu2wHVnk+Y9DW+2gpCPEd9QhG83AAGANy6x14jrkBNHig+uLaxPjjDbZ+Tc
rB2Z63kkQhvF2fDu6fD56VgRt1J2Fwwyp4E9UPBtM8ameRzuzyoc+r6Ze+48rCavfXJyPDolmJtx
QomExUkdnw/gOWjZRPQ0fPkzqp9+3/wWbmei0FfqiD4mZbVPhLYxDodfUORUM4Zl8Z9KN7n71PvT
5TlIWJQWoIr3boqZIWDrieAjc79OSxq/v3Az3Tr4264KjZVRZWZD5pU2XQfMD+MFH0OwG3E1V1rT
Ns3vH3JCnVKj7h1Pmp/h/MRIhTLQD+QwC9CFkm4C85BHQXV5UanxO+sDjNRU5yQOXVaCFNKBnP6o
2TjoFK2OsgbOLWVcFgUIz0l9HHWONP50AfMVdkvAkFAsJ1+H0v+WfIskAzGtfWXHVMbpfjReKhth
bc8G7sEzp1HR/VpQuKXMxEvHZYJSMhjwhDdEFFlGGDU7DMGlXUN8vUG8Luz7Ew/zDILvZahTjLGz
Vet94yeyVT1jDY6t+nCD41vUB86jGm9xm7pjVy9vGXXa7Is3RSlb92oAe0ZspS3JElW7yS/ZoTp9
76WCaRIwdJjvTUx12iy9ZrJLmdr4ufdww162ui8raY1uRkMHvE9AMNk1Hw/WaLyyPBCCjSGFXku/
CyLSJAeVLBuxSO6v1fueyxChnstCM0G1RmD62x/fCjwMqvph6IhTyd97OLukf6EnSxDsx9NIic4H
Px8IMRb2CW1jY2bDAI+ihIda9GgrL9tY4H4M1k2g52Y/f2rWTj5shyYESAV0MLYGCVjDsoialk+S
ixs/YfSFJcpqQ+lxbGMPQd6RVcoVD+810X91USHh6k5vdT2LeIghyvTUHksGlQ2Eq9lvO2hzk4ER
wFOSJaJaaXp5Fl2VxwZ/eDY9SqgDNNqsQ6H0lcN554MOTKh/rC54FNKt79odLVLIJ4g2Us9JfMye
rvrJSTmEuCiJMPbm6ouMjR/Nt0kSNMefKU/WmYDbAVaRRZiE7yZUxCCyHFJe5KUdT+CgaCa5zrl2
9MfcYYZKmnFioIBR2jO7p21vfUEVhklG0vyxZHDBVc553UPNbsFHgHBAdHpTGUH+r+BcL8SP/c+r
q02b/+aMK0xH7eG06rwX0huplfDr+YTS9WpiM9nCRjoAcHiS+rju9gpWCcv9+KyvKDOFeLu4YhiU
8t6SaHWCpjRWpUqWIPLO6krxx5OfeqQZkf25ZT8WH8a18IOUHDA6CDFp3ohg5ZXfk49y/y0qu6Og
6O4knJiUMUe01Qvh5ia2zG9yjeQxdoviisERoR7E8eiqgncICM+tJOhkE4MFeAM2p9cH8l4rue1y
gHCMDCAjsucNuTYeNUNDvLQ0T7x6cwm+5YVvhoTzlORJeqbv51UeqmWDqnkRuLSf3UJDAMisK1qR
+EIZouxOJud4Rq5tB1eafWru3VR/5b8gG7+wNySKBYxKPCEsXMTm6UFzNnLB8mz+P7hzXoGDxwVI
31x/d697VwhV200ob9l1w/W1QQhdiVOU7x9/ID/LT4HkczqkmsFGQv2eiTgh0rRfIA0ozC5MYu08
x1LL/BVu8rqXBSMFJXZrbyk0BP/Qfr+z1JJgZSMY3tOpus+wnaMs1LkptC7+1ED1geXkoBiOgQ1b
sh9gQjpfesqFGxokmZTdgsJyOKfDxokQtP38NjqyBz+DCcMZXnjqBObFxGrpJj5QPkFYomX2EOcN
PYjYIysWBd31x+EQVbBMhIyaW7SmkdPZdrHV6LYkpoNqCDbPqTyDqIO30jHhnzAhJVkx7nOfIQeZ
e4z7tI7b4xnKY7HkdbW/osKvUr5q9FWbTQmrS28YRHKi0BJBNb/GDcfebicUHkD/E/54HH8a9P3q
A5PpnmQQhGUXiie3JG1rsu3hjPh4Qp+EwQPnbF09MsDC6ciWtEsHeAO31bN2J6F4jTL6BesHZJlP
D6/8bl9uXHGqxTITTscUeTnTwJr1R7YCV107lIMdWK/uFF0oe00yOmljpblVwOmkYl7N0CMpzB2G
mGQ/RyEyvtn3N4j7TiEvxf1UVQyiKdY+i5XdwZVEAPg4oxQL5HYfu9h46ptZcGgnp+jpjW3gC7BN
HpmMh+Aybc7750OalHUTAOM/QH5iQ4S75XuphW1ZaXz4A/YNQU9o+7othyDll9MNaHte1FdCA7v1
4Dr9yGBkhIWU4W7EVND5rt+nB8RppOr+ZWRvQbdnD81aBk883Bda4gQSiSHwW/AK2XpesZmlOlRc
eo3fdO9lMq2JAxsuh5bUc0rdyYgPHiBuSiAAz+Fpx5gzRuHBKQAEgUI0soxFru1EvjNiTmZ4nBBD
c9BHD2v+j36tg8wUmC0GvZBdx+zYSb6ersFZKH/qbpJSm4YvRz911tk6V3J+FLECI7guWnCTGju+
0KZJzkibU86bMJbupG6moDLox1STQomWNIbRjquiqjO83YXzzzCAcDZJABk/D7Oq1KNyf+nqtPeQ
h1Irxl9UjxUj79LXqrurThSnJA5qwt78WoqicTkjyAUXB8ZHx7Y4EUdOB5+5pZtZWiIQralW5RO7
BfWpeUUN3A2cc6nBQGVzWsaCWJkqFuAiT6q9iuKXxOPNRUoZ8GNZszrcjJTT9N+9nueewsmuXca1
pwF9tYFl2PqCUkO45wAgRr6MC0jQeHNPkSH6lQrtD3QlA3MQtW+rbwIHH9exWJ95OLLSPKtkvvpP
xCgAjVU2cX704epwzh/jIHHW+SeQBUn+hBQHC5DXL7rWEDN/b/rprxEt/rEGjiy4OvDsO9cDD4F9
zxmB98e57m/EXs+7+9k8nJeOzYkC4P2dTUiKGlmOj6npuP3ulxZ3VuOnX7DJznmQQ4XA9wOekt5g
9LM7VRkzlyadP7s1VFvsocAHIpr08SC8nmZXUozSxCWbHM7ryAcNbPBz4nwFYIJslFLgCS4Bl7z5
7N/vQW3vLdQj07LB0OAfCTtunnwmzZ/aZJ0dllq1XdxOxAtiltCDIhgCTRb9mFCwoNe3BGCAWYwB
jRUltyVHYyg4OkuBRehRD603dQNA7Y05GESyIg+Ikz+xQyVNsiTKtKKkDXueWIo8R5YY7gbELzNH
6bx4uhe+7txcIwrx2MRJ3T9Z7eye3OVq4H+JwmzvzZXW5WtZ+gfb+BTHXdSmwa5/JdCDJshzvxYA
LzxNMmmhZAzdtwbU4VUHM0o4gQ+yd+oFUpYnQR6hW9SaGCbk5QWYfG8pEowfYTL1OzQHMy/gvX94
YbRTQ72P8EN7vj6WQEM5g9G7HVfENWii/Q24voTK91JxRacbzRjCkC4dID+YV+6ArgqpuG/amVga
mRMKoiT7ppHh0jxt+CwBWWygS9Ut/5YqK34Fwm3nqUEM464nzbLEwwCOHfoB9NunPYLgpTtuRTYW
23f0NcyliQ8UqSu5nLhs14Z1S8VT1h0LZUzKmrnk3i7BTV/sKlynRx4nAlYx5kW+A/lRCLah0A8J
JCrIBRRRVp3NuaqcKUZsEM0/jK1j66/KnNS8PwSUtfIt2EhVLyZ8Mf3GRDAjb7ZN2bw4iBPxZfhu
AaPB3dJ/aU9sF1kAkZLXTfUvPH4wnJkhcsn1V9D315Lh4u2NAoN1NWcmH8Z/X/3J9v+WlLx5N4ZI
mLRXjhjwt8bcDXVmLTjM40FUNkwr4tdmHAks9WxFdYQ0/1NCmNopJm6L7MN5/v4zPOkFuFiaiyl2
NM0esDKl2PXwhKwvtVJ6xhQYy1tXIT04vdnuPB34/ES1VCcmR0xcLHPkPOjAM44ENQHtZeyS7a4C
ch53DP0rIOUu6E+v45PBlrTrVFMT7PvtaOrBZeOmclWnA7p+OAIN9emw7QstZ8ucxSfar8k35cl+
cEH99C0D9FHcjNsF3yrygvyEX1484suZ7Rm/F3MsftFj13Z+Nxki04nGq7vrTXwA3PQMTvtuaEpu
EjpKJOxf3A73cVphmk7DPWpKUc93YEd+9KN0SCtrDu2Mymg6ou+ZEXOaAnfdmaTxEGsP5bacfMdQ
/mpNLpDffz3i+aXS8uUFGXze/AhNdNVYd4SZVKCqTFU4XJxyYGwiUpKCXTZPxYDy/tN9fpEocsJ+
tr41SCn3+2lpgwnSX/WZk6hfiAIonHeoZPI8cWYHPOnAH3MDfUhnvpfMJoulELmZxKwcjdxRjC98
cWU9+wT3ySKwEZuq3oZwLZ7vZc4VLbxyjQOF7oKYC8FQBkc5JSz57m1bCn8MAGsaHJK7ntcaPAUl
iQwProElE1QWzMrDVr9lHjia9lSzpQYZq2c681H71kvHtexnEJnOivtIYvESCrp808HtWZHJlBHk
nVmerObnBPv44OtI5vscq3zymOLXtaq6qoHrWH5VWNV8lUi8T/4SznMyYL2f0LX9mJC5ADuDQ6iJ
Ikus2lrdAQi/uO+wLlWtDlXYyYCqgSWrUQ3iXnHA/174PHTBL+Z+bN5Wz2AzlxkLO3DQBhOnoxOt
rVqTxr8AAqUJhS+GjTyzx7Pd65PU+yiYGyFQSt212xi/PqZCg1hJxpyySemL61hO59+fjH5EYBBB
saW1O+tzscm266l2jjmCWByW7SNUNrjOSc6piaLpuIGrRsvvxkI6hfXDNpRVX2+peI1LY19VWHLq
F5jjzWq+8X4wDEMp3zdOcQ9VWXyYNZHD8LZA9GjzAEgRztQw1uSxMgcOLVzpwMnS1jHsJ/eri9af
WQcfg67tN+tPQ6lhWe/9bLAEmPhWfjbybevXP1m07PtBBmkyqMSFDFFDa9aK+KLqspE8MQ6KKKO6
r7CBWbRCvAw733rwffaVb23FqVTkoQoT86LyK3IT5lFyZuSLP1eWtahgBrPfTkTMp2UM3nla6x71
oGfgVZpmtJdq8gfa5jb4woFyZW5+7tkK2KarKEF/L6JM1laXtzcT2eUun2UT3j3kWKbIcSbzUYs9
BiCN47ArD8TCeK6J2AiGB1iCEjnGlC78v+XtkPfEDnV6+nFVDH+21as8JGakY4JHM/9hSpwhnm49
YbfrPEdo3yAxFj8b/nFdAztJo93UHFsXWgG5lf4Bt0fHEgBUXEHTtVDd7H4onMnIousqSkZdodSU
yqyO6fuXMhnYMWV2tWV94P7kV7nUjph7b4+KdAoicpN8b/4BfDd+GY0Fl7QPvCXCyQ3tscQYgir3
jSmSJq0hl0iGiAqyq0GszkzRCSrZ/29skYBDwbrIImDEiHVYfklMsCsXw/sYY88J2LMDlXdFy4Gp
YDoUjQRX1kKlUfUY1PJiKKYs5XUafJ+ZI6z/s5801N7NVJB+e+RBh1gzm/3rqY/HWGIBOhvpipbC
noV2fjSUh/tz4Gn3SG9dd2RyrJyXPVHx/eYP4lWFpP0nF6GVa52BbqAJ7QCX44ELIrXuMkkmCITP
78UDPaFaqy4FJatuHDjLqWoEDj4XAnDk7xDY2g6TY6hKHT62QwhW+HggPz5bNU0cDkrmHvKnGq1h
sK97qiMSYyts6zufa1y4XsM90IPTXox59WGwQEtYrRLfdqwnoCiR3nx6p/WVBqbLqiGRE4ma5FYN
JFjojenZ2XQsxYJGlbGNKErIUD3+h3s05qlAOuC1ZewkyyvEUjptQ0wOZ2r+IKmCz5L5AA4dCjiX
gbBPwlayVjAWaxbdthFQEyN7q9Y2PxzCGIJSXuhWfRpDcTijVjH/IDhtxaV7CUx1cnkO3tEzUDW1
vMHucrh5ymQObAl0haXRIod7WrBBnsbBaGw5p1ywobyDNGwW1nghPsWPQtcoEGAUKmsJp6ILJbmQ
V/jWnCBV23hzV92HLaa+3cS2KOba4RQKgn9+JAkefmGuNWgASo9kT9fAyLk0uAIsUfpRXsbqlGYH
Ura6n0VBLcJPMm7FjOHmwXRX3cO2AxiagGHqVry2a7UekkcXfkvRNsZOu99SLwSvp04M+YoTXoB6
j6jxO8V5OmK7mGBXVsCTyejgioaxKlUTLwnuuLyf1lHYXhtwpUYyUyGq+BdrJk233QOr+HTssHWP
eK2wOOebQQh+kevqr4ZFGWlv4DgdbtYka74UrqkWSk+j6GCJa+gVqCWO+ywaQihWlM4vXuKcK89s
2w3el9QffU7ov9JmNqyS2hcLFjWYL/PMqo9mS9uIDeGQEHyfcOtS+kVp4wBQbj8jVwzMQBLilFIS
0kuXiVAw3cNvAglLzBxRQAzl1mzy35owdkgPaFl4oaORwO9PCDKbWS49QyZA/cfFa4eYjX5OvzHT
v1yqiSroeYe54PzIXMsGp5KJIwToJ4qseB6rINlV7Fe3+G6Wz0/TzJz7PXaeFJcFBN7b1JUO3ckN
od2qHZj2BUzXxDJiBeltc0/n4jWFKlNEfR3cZ+OpdsyVPRqDWlewAwD7gl/PYiKikY3WDLj9967p
kGaesrI1arN1OYdX3Cbodhs/Dd3hxop1/8WrJka1ZzAk3jTSds0BTyWGV51v9cNG3oxoja3lRb1n
4kjNvwF1xfDsiWcC3U+P8AEyL7VwxTIjjTF+2hyTgWHsjE7Cj9GNPC5OOXKhq60fcB5Xuh2+cMgI
wmKkVCtjwbXALMHz9XaHcT25+KGTvgu0j8BiJKZTrB0W86UAkY2hBGU4fvP5KSJ6JXGLvf9cKHRj
iEOjkOU1EHmrmKnBKWL6halZbMGRH0MUF6B7hLLDvox4nKmuC7upRvxU/O3RERRx9N1Y2NzD2vd3
2jLu11ytgZKryc2oywRv72x854UcZ2YIHVDkdjXBf91FSqNN9/GBvrDUKYujrchuVxhqBN6RQU4i
/lkdYYN9pyAi4o1qDPBPVpfHJmZeOPCU5CHB62m4Qn8eEEampYCCNvwCRC6enDuN1oaH8B3MIxVf
YIhgSJaJhImxuAKs9Pjs6YTktwaYxhK9WLlgwgRqgJso1F8OnsaI9b1rd6h4r9kmbS8w3QCqWc2L
EUqpmMEU4qtDRhBotBaYasByIHOTaNEZvftiwHF4MzM2GR2JiqgNT7fL5/VALSSU3UeV0FPP2s0v
mict0fmY1AWgbeuWOcYp89Z6nB+q5BvtXV/jEag7PQf6GS2W9FeNrQ6QGX/t9HBtnaiESrD35u8w
TcFn08SFEWYcIwKhDfbZnRztrxBMVzJYD0IkBga5uv4zuLSAYkfy0TY1nvwX4ESgTFr3ex8UHiOl
Blwi5cRlLg3JHmJ0prCFIx1Y5T2D+XzacdXrtoFcvJYzq1be8CGuiTXVNpLhtAoEzU6kq0G+im43
9a8TxvUzCbmBsxCVZBL7J3QLztmJmc7ZUB+bujGuFul0+OtOHT8WTRzeaXbBlF2lG5no/7sPYHoL
nrG8rNxpaGGUb5+Bs3qaEo3Nz7ileCfhGCBWkm3Dc33AlTEFMXaheGZEcU6M9c/7AWmaYhuhm9l7
g6LiNFfYnqB7AiKIvfaFpm4GOTl9z0GtA5ta4m6UV2oiiDM0dPZmfqj4k3HVDYkmey7+kWNlwCkO
toZJwU7iT7IZFuO5uqrvrYIXebqsGjN5zVdST1cCZdWn5xK6gJYDb0X6q2iE3dFHy9lVRw0qmUxX
HEFFZgLY3MV9bv71aLKO5BTOEtVrNT5U35SOow1IdhP52qtFSv07qcu8dK0MdT6dUKiYnjY9u2YH
O/2QrxE2SPcOZ6shkous5I2nRts8R/RqVtNrpdVZ6A8Nl7MeH1MvCWvm5ypC1bDV3jpUMVc8+zhT
doRM8IroXpobVw/yHRfPqMTjIb1EtqfqLJet6fJQ59aTESvan/k9PjXD1TEYh784YtiMQbQlYAhO
mgBTmJZlHDxXOr/CmPDnn6hOc9R2FQJBxx1Hx6GII5D8m/AOmB1PL1a+NtnUAvcfCb9qf4SvAjJt
73pCgHIwWtV/Jc8rETH5kbXbpnxFlXCPmbsIXNiCcV/u60Mo1xIBv/N1RvP6w8rayoUI7uGJ4Yir
AxyADtjVqsDoJWUDC5G0PY2Xi6cfV9wdrzJneMRbErpq8NPYtEB9kU47I1mTGk3M5HVYGhpp/bQ7
Ks2SboogCs1nj312f0FNH9JyxN/5J56zW6gQsmDq+5cniq/XlV7pu5h+2szRjq5JMaqktk+1uiUV
FxFGKjcaZsTgVSSbm2R11Vi7XTARh8Oe7GtuRLh0BqumXHrNczOPbl8s0lkxiMCzKcRWh4exqyx/
U5FPdlNkH2leQRE7k9zBlRMToUgN+OnZlwIxo+pRduiHykmEdUbfQT8g4TWN3ko6oBFbeZOSE0/k
iXNB+1srhP8/g/+JcpWZovuZQkF+xlWTjvaHTHgrTZa83qMkpiLWO3qAJ/Z32SdVH9VLwsEC+Ins
FRWOa6KfAw6eS9GTyNX5Ylvg1iujwjMsA9+IhZzvUd87GTJdovHP2y+H/z4xefIa5CrDMZv//fbR
l13leILySz93XBsSsBFVvicC2xK1joEfLRpvdvaweI/5WM6n8Azx0wFg3Po5f9kw9ntD1J6M2Njh
qbMmtFrzXcqYryPX2KXjeJI/UES9dChzwqR72LEDvC1Srewpa4nuYrkhCuqfIHZ2af/8J3borEYv
BBzPp+rlxpATavrgKyeljzbZuijhAOccaA8LbsB5bQm3DNf1jAUIP/nxF7UyEE3ODCG0/Ei9k3hj
pqDzMMJgcefNnvccNBan4gd1/8LYs/2k7G1onVMWYfL42YMFvdbHJr5KtqtVuGSCVPjsga6LrSUD
uGwlR3K8m9vwpA/LUk+MBII1XbR2myFZydcodemSvokL9o2i7z9/mTgZOKW9/P+YDBavjNUYPtou
nwQlQB+rtn+8F+wZVelNzTeHMy+7Pjq7vWoSiN7iRFbOKCqcuM/PS4yLZ2M8GelUo+7k0Frt3tct
QES+sHd3m8vu6t+l0EKewO4y1aDid9L5H2RrHKcJITR2z9eBpBm3Ctctvv/c34Ebf8zKWbG+GnKY
5vlTv3IS7Ul7PbnfWCuQ4Gw3ujDydzoRR7jATYsnpI1zo0cXrU35z/skCYud84J2ZZDYtyCA5Aiv
lQICNybQe8uO+yYrp3Ab9RnDP1ykEEPu2eIYWzLzYW6F9mJiYRvwXwwQ3kS5qP9KllQ+dI5k9cwD
3Q3Qu6C9TK8dyKcHhGHIIzrMCfkd4mmkI4XotU2aQFTlfmwWbExyvVNI5hnVubY0LqBa65HTjhSs
hQuwmOFHa4QnslpJ2Usk1qlFrGtl6xwVQ2o1qf9XdZmZsCPzyF1FIdOpWngQoNfieekh9h6RFmte
I5/A3keutwbAgAnTVmxZUIGNT36sdvO5VvcePVxjYi0GS/hFqDYHDHJpybTJYYOgzO328EZWuGbi
JlA4S7AdDGONec1cUQlipKEbn/nCHsZoFTDwGSyelgq5pPWUf1hwJYS/2T5xcSLMHu9OVtmTqw4x
w2Kicti2DZU45WgiHKPCkvASUIpoa7DybzXQdFZDe0XdWcOHPPBSAI6cJoZvvlxKjpzC97OnQ7xm
ydpxEklpeAeGp3rwgQvz3KOH9eM5W/DpUbEiZS+f3WENnPMPJNErpFyjh2wvYQv/RuMCyjuUJ63u
GHusTZiEPk61jE9e08u+6jgBRPXhwhImagcGXyssy7+svQNbnZiO//3dGnJtbbtl9iiJBUmpMA71
R431LtL0Its4zdDLPqUDg3wn+41HURaxNiVmNF4m8f5rhRlG0OqWdOz4T6N/BSDEPbD0TFpUQg+w
kCCPdl21/gGXc3A/BRfkV/wEHXRgByFB+YiOCpIrja3eAG+qImTRTsgwk5PEic+Gtnev36e4RThO
3XmwBncjXZSfvJLLoiijKeTl5HBsvgDeKfx7Gvw+vON70z7Sav5QDsVYAoYzSz29P7ftsGxmYA0Z
83K8ltxIlI20fgJIyYeYi9LQxVNuBJ6ht41y7fCjEuxZ8R7OTsXlWaTeJ+k+1rssVOsvrqfNbfZy
esEQhcLwowdvlKsINafWpNuESRUcw47Ea/mwuK37pf76eqWRwBrWZz0XLwLoRox0BvV8Y8cOl2iq
jiMoRuBNlVgtR5o5xM7ob9guLRqaqAakggbAn20hNjP/yrtZtcBCZduzxbZTUGd+pWy7aHOw9rbu
igzNprsK43YD8+pUKiOkGZEWuP5IX2ZuZ7tgS1TgGA2v6XXTJIOdOdfDT5pVZHW8+JDa/b6fUXvv
Tt9w4Gvg1HKxw1EzrxqOZaZ6x719zeyVIzBbvGKJRjfQUqVquKebS+1HNbdebgcN3C3A2V/l7InY
2zrjo5j33h7EzsX7biHuKL3pFFC1Tuyu0jjE8+i9L9opyveiJr5Sft7OaIJ8OG3qpC1osZPwKH8Q
JQCEL9xhxP17WIXBVpD+9u5ePQk6ghcze7YYvj6i7ce2BS/pbmZVYZUMK28+ejEJVx2tRk0foKRm
GZIF9m/upKhX7OZV+KvWCkEgH7MhBfgDx1/zkGh1K8XVL6/b3uz17TRdeFPLOYQsKU3JPwc7M77h
UGuLeQTpK6H7kqFzEVMlOBdcHcAv3wZbhSxKE99t0Wh5yd1SHqq5zyEiAR+LfjALAIhdwdaDRLgS
pJVBLw6K7OqfCGwOB15Fr1be5zrMurXIwKvMdJbdZggzaCNQzMLAl6NiXiTTLltaLAirCXDGcUtu
m/hxBWLJWWPqPM2ZOkiekYMgjeoLRa5maHCl3ifHCpBNCHhu3mvFH79AHBmxYqXAOOtZtFirmsAK
80ehHKyo1KGZwRhAGpOUKBHsS8qu26ZvN2ZN4PNITOBYXRV4zsoRoK28lzosP4Ik1BhIwRGFpAWL
0DxcgKAs99gZk5U16abagT9n9gXLaT4gBX89oPRkhOqFrjrDFjrG8L3KyBut5VfuLdMm0/Ejk5S2
ZbxwZyVmqY+i5OLNgXmgjnPEFyyYkuNDZZ+7PylcU319VbKCBTiu3NBgiaJpTIdXFldOWvHZ+eg6
svkEEcld8NktgX4iWpZP2iRb6JXrKqrKwK5xUEKRQIaAepw4KyoI3HJwxLBfrHI8BVkNeG/MBtVl
+UC/zTn3Zjzq6vixYmJRAUImY168sRlFGa9HQwJX2/gmjLONBkLA5PXYhHfKOXU+VOLKiB8QTHph
hC5r/hL1/J4cpdmiDvn787DlfPRtr8FzbhxdzGAJAwvuHSDtJHpBe2/vyA5G4IhxCNlivvkDMqU7
4PX7hIZ/crd4d3EFItVw66pa42NVkROKmvSPBHAHyMeK24j5eRXwdL+rG1iTUEvZJrIpBY8QTGBD
r30F0wHa6zyVe9gL6pthkC7vaMkNWwVgJlB9Z0l7NJfu0Us87Ue2XFMw4HehnShOa8Rx+9mo5Kr3
8igC/y/Dlv1v50waL/nmAg3sJLoIbTvRjMlkAXWRgs4Zm1XWA99wkeyjRz7es4kQPAY8BG251Xam
jkmtacSFJU9A6bve5jMQ4t4ZdVsAeljYsMv69/86XL89/gUBhTk7TsuUDyeIaRIx6i2rF0rdA7PO
YePRDMlykyJDQE/wbH4PPxKfujKrPNTL4FPZSUbQFGJwblDDHdWEQH74vTUV8/vW6310saoL3pOD
cLP0d0BpbuYOuVl9Xm8jMb4E+g6BvYpDn04hf3ZHlt5xcffX/GAEnVoSwG7dMZP0/yheBQ+k6ClU
0e+7KKUBgDg0geunvHnSkuRgU7Q6XVi/FwlN0HSiUZ2zQWyi9mHi1UyMlIqj0inXvtZgkH+ZwUhS
naURjv4ywI7PqjCcQvRYpdUQJSMi2ujGSm4tgHV/tTiT+etExyGsKON4j5jvcp6IJUes7rZ+LyHw
bxMzlVSYqTH9hCLyriIPYLMxb9lqCY7A6UZ+8gC0nEesQtV8ysqqFdSd0eZrnZK12WLgv+Lsaw6D
WqNmWrCARZd6XhnfDOhCwBpqwFW6Y+MJo4PK+kHWk6KMIKUAXjUzSYuYgtu+nBKKSp/EgBSo9c0q
c6Hu/ot7EwRaC/NSsPIWEwPQJ56rsK3KkPoIAAnpzfreIVYYWHeqaVJiVKkZwI7KpKwsr+Q/gOBH
i/+1Gvd/pSHl6AD2wCi3rNVr15Ue2iTm1lt73sZoNKDIraPisdzT+y22oPFDV7TxkopLNZ0cdzFf
aRxFA2KhYTA28xRzCMpA3zh3JaMOlp3K7Lgo5rJuBa/YDJuRnn5THsrcGszz3T3eVw3Vtn5bxcei
MkC1Qz8JlcUJsPzGMpbpVk4zlK5vUBSt3AICfPuG6RXvvXGhXsz/yhOYij4/g52qlJ1uo8QdvjMp
rdqBeB8MsbBtKQrexrddP99jYudn+/r2qy09S4szGS9YiUpEizBu5VNmOD0+IS0okDQYFSQ28H2h
HTgZnNcQochE4mDPNznACQgRJIY9wX0C9W1690appqkwDmGrahILCNei612rY8Lo5tKcSMmF6fE6
XyxEEGmmys7bJPWY4FpUWdx1ot8z2A6O9URrrdzLktLpWDVvQ6Lu/5KQki310Ez4jK/NFCYRhDYo
rjkEw2T1Ppzay5ybLamFE4tMCbicoI936bqU9GoozDIjZ1dTmNuzkg9m8H8z41VSNH10CHP1z11G
byGHSTwd6TCt7dOJ0SPw+yLVQSw7STDhv4bQxFkS7LM3PIkAGnloa7tTDNiobMJegFS6V1Vz5YNg
6hOrmuO5Ku9r6REpgxI05GHMhk+Qer896sF34qx8f+nYDPwUBwX/F1CdO8OUOiZHklSBGAmoeDxM
4i7ozZ3izmnA5ahJSHLna3OfTgxEzIilBKCQfdv7bsmX8sxmgmrA/7Yh3cIm/GpADhCckpjUlo8M
aYT02GWRlcLoG+j8w6iGP6njpQ4gksOJ7MFhtMDHkE3WPE3ARrqg1hiNbph+2zXr6GYBvP3JBSEM
Wz/KVoH+mxbi198xOKnJQV7nNhT7pnETWnihmKhhpbwiR0K+XsVGuNqZHFZnzNcPX3G4CgH0yKnu
hVfzRzefTyX19kjhovABsgfX5n235/n50sAH56WvHyCenbSbRkOXUD2sQnZlxrXsJQGzN5FumsJ2
pIqxsgkl7vfbC55ODX0t/35dfzq5uhtR7Na2NljVLzPcI+SmvZAzWliciZhWjyNbp3NkrC/J9wjf
5ALgxj/UMYWfX4nQrEI8FWAt7P7nWaG92D7B/hRO+FAwnNui+JvdbmKnl49DLP96LPw3iiSw+c9+
vAKp8gdy3ZxVwTAs6LispagpEW1bcDoi2qtWQkb9vsoP5RQUgi+IBBL//g2f/XyUUeA0eoXHdPJR
Yi9LcBzx7jDWfe8KITjbzKDBToqQL1iK6n5lFWfL0ZlzJCqlHRgbhtQS/EF3ntvdf98y87XBEgeN
DKe3X18pdjgxJDZxld2L5Wi5RvvobyD/Mn880ViRmq4hU0p9/7Ao1qbTpQYkvyNZsgJcxB3LyOT5
3+JCpS2O8qBcu0V8DDGHk6CbtY5aD0UjnxHeTgALb2W6sOL6H6DAeEn6GxHYk8SiGHw/6lMLtDpT
u6QMrRvok7OwvEtKSCmbUdcaUK5f6zhAcf7+hefmJ0Nzs4QHwy0i0Xts5KWVY77qOR6dTz0rH+MA
zp1SPg+1go6o8NlH4VIv6avkoFbtvclPwEr2d4V+uBccTz3HNVRyqHwGldFQczC+3IC/4DKNC3Mj
qAMzjzzLaGLmN0uakkT/D6lqt1JiWbRRWHek4LWfKN7r/XCX9mXiplsH8K7fnuungd5F0bKjeiGV
jFeKo0uZlk0UFexuVEfJf6QiyQ84QlZZU3ZdfKMTkq66oc8Ah2rLRl/1knCHnRN6jfnQhL5JJheP
K13LSYqE47ZflvvJSpNrGZXlOasXNIXj9sRrvorrvmAp/WTul3xqw1zZ9/wt9BeudUUduWujRwEE
0bd2ZvOIv6LwWA6AK64EE34Fqwhl+bGQ96eo/hG/3OXvH+jWFUSU2WYsUgWYMdC6pvtY1rNcb5Kp
zDSG24T5LnlDjjCfJRqso7KDJBGNFMiLjZFbqsrbFBpDSUwCb94SHRxW64CnMpGnoLCbjgYaKa71
WG6Jjr1BUpsDXpd3ACTpDqdhzSvXXQnJHoQkB9Gbh5cFqZ5Y+i+LkV4SSboSS0QK0/L4YPbNXS1M
NySZ+2r0RBOoDOIditPRKXG0wEoGZr0Qy2w5sRiP6/joEPmse6TatCmQoKAH3UzWe3DiJlTLFDu0
OZpszytSu4/lDeg10tdy5FY5TtOLpTKjqbwv799HMBQE0CRCH2Ek3Y1V+ZMWdLaarG0puJ/gni8T
EwjsqkuGuB1XLGF34wdAYHrrsogN6PPeSc+r1BibVPSJUTJnHIoqLw9KCymy5YrC7J+4SB4v/hBe
T4LNs0Y5uNH8VIkjzYD1U6TAcLo+RMOhM+PPj0C+AAoHRY1U+IKJxGdF9WLsyf2wIDb7oJITHYOP
16+NkzpyMRbR6mMyKtJgp1kQ/4dGIKE9o/01E/MEuo6ixaVJC4PO1KJND2gp51Wj+v8WO4JWXcaw
ROcuNFnRSsLmuFK8NV+E3mgO7kIkQPWbt4AoGtYZphBCQ94sBr8ZvT/ScmauDEFhP9xigqZNsEzE
XXJ17FJ2gLG4XyFd7T+u5/8jVcZ6T8tB3QFw/r6APgSpNfdDQND6vUy8EACp4mGm+ia+n8vIsUMT
yzhc2q5y7qgbms1lQRZN5G4XRVj635imk7fv7Jt517BbN/ctrZvxwAoICwkjQk1sGpyDDDZLhC5Y
OkkBvYBWJAZUaNKNbEQFvFUznHZ3todFza96A+xw4s10znHFL0DAje9utK3v1w005evLbOv3tCsN
66XhKndR1aR43iKy7/ftHYUAN3pEkZlohaUXwpTxhEjhW3gAOxRgdGdHCP8lVXRbq3dT+V6fZtuh
9xCpANug3DzGPxgG2lePZBR8niAcU296JJZieuPh1Awu5OckHhZcCozadJ4Ygq/mLZTAilXnFJY6
bFduN9kEWaPLujrkINNvIcQA1TMZLniTFVT4jtNZcRc1gBcFr+TTPsyjN7OySDsoFCqeJukpQpNs
Deq606G8kXHy3U0WyQOMNFUFFJ+mNsUPPhyhNptbiB+uXr/PGvIonXDuS4Zc3L/yo7pquQnhc+N2
vVG4B3P6wHvMrqbdoMgJ5gYZuNk7l5xFh1Wcfm33pQNCbyHgbopgEl4l/9BvY+/us7MryehKP4BR
ayTbL8Uo9HolZ+/VRvjg357IgS9nNh6AHNiZP7vPdmHuWAkBJh04SE27lyMKueqSJxQHnvxq/9G9
rCPNCQDyPERy9zhIE/v3PB1jcO4TjaPMvfK2H9XWlChgKEh+4jAnLkQT8Cru9+uRJSceWK1145lS
R2zgfeeNJ03hwGtDpHbmGpKvblom8FLFsPnDPNt/lSAhuoPIyQ02BFBEj/WbvemG1lEobozWcsKs
hO1ekHH7/J2bUvuAjiVshd9YB7fSEfiWXKO8LA8HK9qmhj5jdq9I60iAyOSvStOn3uCWuccFM62C
NrDbldxp8fcBl4hKHaCqZM+aMjGqY7vL8RO9qf6IbL0Qi8i4RTlwuUta2a7RrLo+0ftWc3mzzIcx
IujObgUeB1q2tOywy6jcQAAc6LsUQRI4qpussvReRJOM228Xgk03I7kv9x8B8EWhJ618kavn6NrJ
sV9JXQ7P6zALOPXGt/lolA8BvH72ALQ3i0EQUmpaLL1nAZhlDNsNMSS1LLNeqTnwGZ7ghPnuFDkc
QCpkBBcW0y9p0DXn7ALoigAdXDvVHX/1WkMGAiAFNe44MGe37G0mmjpKTe2quXhzCWe6/LhuvygP
nhEtO+MlwcO3jUrtIfhR5xYgKLMRI3h0+r9DTh6xwd6DYCw3PWJtqW47hBEVmpBh0XVaf8+EXm81
Z/sozNfwttV3y7Jpoa+eLIhv44sDtEObRx/eDmmZ85K4u8+fgJPkjnE1WcvAGAvqWom09QtQcIz4
iMb5hH2P5XcQFJ1/4/xVwswoJee8ZFIzSF+UHJofnv5sFmgktIV+EFeykFFmOlHU6j8RFZ3Ti4t4
Yj9BP1ZTWmzxsyKxb5m/Cwzrpzh3MepOiaW/zjcBB7E+oz027txMT5lKmMW39r6sP4a52/tqO0So
vQWJ7c3pOzjA2M2MkEYltypmotlht4QejNHEnpNvZzsiLGpe8fanuxBaTUPVlyk3amnPB1T4zjeU
5Pc99ao/rtRP1Sh9ZSmnfhtq01P2nSz4l2n5Yb0ZR/8xzlAiqGRVjpRjKbCVK1Oy2W0NcxBP8fjI
qaym5aehRMCo2nxlpAoSUPNpFT1M4tWkAVuWYIA5+dw9Uy1uF1N1CaOjRLbR6o5LaWpoi6Ry/XWr
2i5YoSFgAWNGEiz92ipe7CR3PEZHf8vURjYZ2Ov5BsOIrxwCIWeLL737YW4rppopyBdILJwBw1AI
j3G5V3+zfW7IcsRkEMz9mEcivlGVB2QDlg9Y3i8h++oX4bu6nDBu7MktHYRTRUmbnHlTWUpK8gWs
2wYDIJG54Wa4OBwpWBvePXN6ndRSrZuYFGTr2lb3/pGxZtEmGzSfxLlCLdQkyKk+XUkYH1K0y71o
e13r2haR1i+eSujv9D/tTDNn5xgJiLESis3CNqRQTR0YBUk7iQgpoz0IEsNSsGGudpjBNXqyijcA
rZLesvRa5zQ9GuDxF/rv/hV5O9dIilPum5Al7qYrEtBzksBrr3loOuoBjXOvJQwxerZtQwwMUpmp
1cAMQCg2l3vkBOagCH1qC3bGLXcmo3EJSqrALGLXwPnlU6LpdeUsKtVHlZmbuZ21S4RffgjfenzD
aHrjG1FkG95hb+Lb/cjow6edcUmDbUFNATSTrJ1W3oT1zea5AY97Pt6Jq5O6mqHaYg2mINeOBKYI
/642OSIC7t/kjHlZtgtdXlnCbQLjPuwEaXYIxMp4sIFt55s7HmhMG5fSStgUPYAMJFOw3f4NIbJD
6P3ES33heiAUhi+Pjif3yOHip2jlaP3Cfe1GKVPkWHldzaWu7Tvk23qn4aJKONnf6Lp1u5e4nHNP
MyFghJL7tOVPRNrLTFGsk2gaSk4QdLPtGqT664pJM4IGDon/MqM7tNKAdyKNeV5Rlf31HsRkz3+l
4vmjYluBnz946kKOPPD4PWyBEVYtIaNxBHPoQK1PTmKjDikXk1tx+X9wDu1jiqTtWpm1vEsmooLN
Hd7ApJRgbsH+q1sKgTXz4AiFbPq3eiTiahBA26qPaL7ZokuWC1OahKi2ndgjw1Yv2KswHODyutFf
FcpITWt1rI3SGgxaTXffPELklvl9WajQjTuyArUC7lJjflkd/CITJJZNjsitsbRCxjfARD66ReMv
VliRuiBThWGGSY682JIcC++otpxHiBA6LFaxjqFSylu4gVt5ag9hF4xXqVfqk9NiKUyx2Q7HcoUh
uRAceiLHf2dh3i8DiKrhvq0tuFKHmtd/zrrQFXmzzyq0LDVfi5KoBx+thcSg60HlvxMeW/DMZOyv
lR07mV6U6jMw4e8p21ReWGPplhc1gsU1VVQ4/9/hqqhCCgdQwWSugdr5fvHB8RLIfxftlucckWiN
4CM+sTe7ANBKvEEyZieqGF72tkO62+iODzVaPErROBP2ThqDoYVfKeall1/8p8GjuuJjTc3DUrph
We5WEoep0fvIRtlN/UFYEVyZ1SR+Ugs7owORvnv1EaGmyuSWNKoBvuWiCsxxy1jNFXxKljz5woMC
xh/w8hCqMgU0LCURj2J/nW4fzh10sQovh0kvNUEaVOThlDN9UoZ5p+9/A7I9+soEX+bji83eTir/
39rpqc33p8ICEowf7pd3cmPs9KRk7SYeMNJHBGmpa8hY7S2uUJWZqGRmxlQ8JwklqHyuiD6z5jpg
sDv36fQC8c8vczAXv6ZfhtQvGos1d9IDEPGJIWQJU3tJUXt64zajCBaG/jPd4BVK0HUSRS+CN4ka
dsNruBfu+ifxDauTHJBXUzjzobGtPzumChF5rpTfovAji7N5JzXJsARKt5FaTbtKyvpxwq6oDJx7
yfP5QC7snAO5TwyEUO72ZoT8mRk6J75KGQ1G/kYHVcsCmqr7liNAuUBc8eBz/6zEf2HUm2S+iouA
ReIIovWWU3bGXfJgldmlzSIGvN9+mU3eM8YnLx2CVRk7xQ+yGhwL3dcL2N6AytFkUydJ7vnw7RYU
GtcJZpObtnOMU9xp+sX7uZ7cB2GuGVnbnhmWIn8hpAQxFaQXOHrySoCExNcYk3OFQZ+wyj6eWvOW
tNsNfdqmrhZTmGOsg3tk1RN9K2dMoGo6hr6T7uHs1YUNm75rMROiKH8qxrzl+AMURLv5xqekSAPE
B3LHvA8wcmzVmnivtnPgKw+yYCemdi5xpjzvOeaFfbDHt+j8zbr18lj6YeJoe0uvIys7ZAkSUbXx
XjWn50XJZtIYumVOU8urtfLIYQIhT7N01JkRqj1JV+m3dhvwY2aRJhB6wDeX2AoVEHbZSfqo7+ZE
Cn0k+0mAa+tcO/0KJCBFldiWyaRxH2M0WhxDV85WfiiLX7b5czd+aKav/epwh0nZtV/lHsWWLYCk
vzQjOtEiSxEKbZ1V2Ch45wK+HZ+QB2dWolIFZOE3/eNrU2j4uxs58nU2L/gdC2Hhfcp3yxq+ehSe
cZ2xuAsS828hAuGD4Q3PgVYi33GyuUvUqxr3HXX72Tqsl6hp79UcNRihVpbgvhSJ4DEMCO/LMy+3
g4Go1RMqKG5ZaoBcWZwShFyPtngS0XpCfNRJXjiqTYmWyoVCONcrqHisAnRE1Ljvfght62ZAgZKj
pMf1hscDVtIymbN0aZJUhg5c24GP2ZEnn23V39JZdDzfr7R+bG1z1rc/gpmgQc6Y4A4b9xFJ9HSx
Hbyc9UX/fKyCVNgOxFCtVTVKGAeq8SWAaDGCKcmNE9hPuPDqi1Tp4fD00sgqkqBvqdTj2kdPXtdM
nWe7xf4hrhVb+zyUn+kJZrpxBjOrvMUDDG5ITWHHET4JowA6kz7O2VCDcljsbuLCLS0JpcDhvEnd
bDRdcmM5wlXoOHjmV8zeP9CQY1i5QuwvTZum83dsOS8KW/mTDqDphwBGlv6h+3vpsLG4Miu15CoW
t210EqTLleGmm4uG1JJHlKexmWQGTAjk8tFWCcKt17dvnl9UDb26AbaOgm1+3v343RKYx38m33z3
Z7o/5m3anwKN1pVfokEkI7Q/8purd7UFnrQJqDum5uN5yEDysCPH1CiC0RbO2Wds+GzUBrKM3DxS
+Y2Pprb0x2TjqUnuXjryvt8PGeCeQINby5xA39JrvGJeGCsJO6U3ZwHVnW/QO5XnfjKlBibP1U07
yt3BPr60iqkWeZjyLWr3Mdg9Uwiq4AVyk7uUN/dKohsJdYAcYNcyArY7y9DePQ50FF7TqBMeAXVD
KDmhu7OvQ0liZeuvokAfwlf3TJU5BLnPFALSrynWRfgiRIMhO+t3FiGo2HU3/BbH9Qrr4DQkikUt
wFO1n4MAhzRoOKNUHGhjZ2QKUWNEtyjNDYoRik40W2ff2Kw7ODZv5QC+AuUYTAmgBoEHEgoWdwxN
DdiitSj1o4esllpscYW01ExJes1BugO1O5kUixyaOtipO10a1pgd0jyzI8K21tN0OS76glQDOg1s
T1kQUg+/i5gjC6CF7+0omquaPod4wbACFaFLMXQi9wATR4e0Vu+ybZWT3BAceKJaP47FFrTtDr/g
EIig+kVvQBYiSfddDlfpZX1N67+Kq+ZKjE+mhHzsdnokIBiMRbcPWKc2bvk9Zamh9+I5rTaMcSic
sAC0345JNTJ2acoVcGLu3eOW40u3HqVUrYFtwx8X4ngYhEmOChHfGwSGMeKKF8r8qNt7IGQ+L7ex
Eo/S6xm7tKfagPQd5zf7tKo4rJEC1AsgPl87uB8UiGelzXW+DA5pZlQEBhTav4mckrNlfql3+Hy0
8AdTfD8hCmnM3hL8slDSAxbaL5pc3yPJrYRuEUok/BU4Oow0z4yztxJxFkyByQ5HkJWPOkVQD5fO
fOwpQoYoNj6bhioBHa5FCYXs2hcqQ6uxwYj3nHKrvQoYRJs3Rs6fVaydvEQd9reDg6nSJkcgUAUU
8sYJIi8khXhSAeR0Q4ZPeTBRf0hbNKxCylDJ+bMJlEpEkaaQYT61BZ3bq+kDPdf4A33gUe3KTUgr
X3z01sJmv4PT5Twd77mMcxZmCBbcTCIZOaLgIZu0AabY6/gp+JuChjcbFivg7LUzZh/FbczJP1he
W4uhqRVRgqRb8qtHD//mY4C85j8B9lRVQJL3O52WR6bkP2G0Ykho2P0/aaVBh+1laibxwvmXXZe2
K+QSY1gobqsDKB9fGl46Hd9Q9XgoR6agkqIcKk6g3+ffTFfei7xNfnxGkCAEMbTDKgJ6P0RbP43l
3Bpk17JewhyTRa4YJmivIh6H3CZKnxxskV4gsho6ktsqYhxrEEpFWLA/ad0fS8zrk0SngM8LsKnA
cTLlmBDRYTQPd+s8/EH8xbR+NEooUdDOx+Q3Ygcz+bnREO7G12BX90fEuVNWa2XeK6fTU2sdDCcl
B2wWlPKfCQ3JHZ1xSv1JBdmG2kE//4Te/QzOf7jqh/Arhez4cLW0t32YUs4jMC3FtKf4nluB1Aum
6yWXaibWmqfvXsD2tEpfaWKrrX7nExM6C5lD1E0KPGczEhmpLdEVGw4jn8yni3V9YCUQICK5zqx1
wo8I52+X6piIR5PW+wenSfCMRscQQaTn08Ozc0DbPJJJRQRSj2FF21x+VOSjXSZix3Kr8LBvmCUj
nAnUz66oPv5EmaPjGK3P5cG4pa+0TCXTgFAlHgTlR4ioOX34ansqgZ31rsNq0Cg627aKlGSdWf79
Wq6iMHsl+vAb2DZu4p5T7s6h0Gf+HQJRrNsbmlzpgjslcoxgfX99aG1MnMdUSpROl2J8yS03ER51
lk2Ody75Qm8pmz4sD6xdS3wUfgm3PIluGPHj1RRe9c+rnWltBqTmfUSx0SRmwukqsKTnhoh7vvf0
K9m7seM2EW6HZe9Q8W1YRVnyA0MmDHVN8dAAZMoNNeuJIQRbM9rTYd87hC5dlHeuA8wAj2MAxQNQ
1NBYasw3LYlHJ/vs7KtUn9jK0Bsl64JDrRwKOU5hhIXGNSUotByXCbBZDUh5OJJCDZvv2SILXKiE
AKpsJN9z/XNU/IJZdwhU3bWVLFiKod0fU1lSvP2zA37Pw1flvePBstBN28QyLHI/Vl5qTQbkicvt
pFyQ2kpDN2P6inO4Jymqi3grgkZcnvxaxEs7054M26aqYwq8pyEK7fc2oKHOyExJXKUCFOwwOT2t
RloJ+hoV69HgQiSHywQCF6owAQ56rBMEk+DwEfxO7FGFJ1i6khbkDnrWYxjNx86GkWTpfjwwgt1A
rt1NQljXSny2mgI8sNRPmvFR5S2PibIcwz70B/crNYHe1L6rKnPvPEUcRwIf0kD4Vll305GALH/k
yuOvWM/px7cq+cm1FYQ5G72GcJO6t7EZnX0e1Tq35pe/sn+8zr6+tqgyw3BNt/I23Z12xttZUXva
cc52LV9FZ8Gk736MrLpo8PnlGCBy27xnQkJMA1A/GOnOrGZ33ZZzo+4xwlo1UzFn9KoEDuG4iWX2
/Z1OrvLOm+ej4yugsh6HclnONHqeq/bAXB4w7mHBckQhF+NUBu10T9uS6lxp1h8mjsU15OE4UhES
dEoLoRbLY6NcXExs5LPiDs9qOTG3NZOG6QxLST2UL7Nv5zexSfmR8lVMA9VxmaNh/W1r1V8TcpQZ
jE4tG9ReaDHl+go0gve7adfu1aEAdSPFKvVAuKNkY4m74APH3mu15DrX9LOFzL+1DnwsiDPPFyzy
Wn+gjHhrw92vaPUcbi2ODrNMk5mfbJOwz6oVpKRBdVoS27dqr4lhvIvazGWD5zJg4343jhbHjKNG
jrE6CxOhPKR5AmPzwMD0W6iFo5NpzPUKdvMZwFgheTG/hYpkK6onP8xH2y42x4M/6a4b3ozt4uZO
kddy3psqJ/w6TmTwe/4wcJPq7MVZyCDk/Ap1CsCz/Kqu2cG9JEviYDq/s3CsH5U6jpbzHPXyoLk0
cTP4cCTpCh76bER0LYYVDlyNqPMcOb2jM6D0qrI4qY4xZn63eF6Wx2+7/4A/A/+rHs/OXToq8xC5
D22XyZVSfVJiTE1lI0anc4tsWX/aOhCvYJAXSHk7y3MNzpG2IGqDPslXx6QcFlUV45XhjayGsBEd
uGA3eJwt5oKB4H3f4wKw1rC+o2TmEy1rbOLOrmDKAtOhF6SU0rdLK8lYa+JK7AiUwQn6QNm3yvxi
zjt7+vzvtoB0mxIYbXR3U2RRi/sjo7e7dV1Pks/10rnfOXW/49nNWxD/cLunnvYXex/524RljTG/
cb3Tb8BN7L89SPqEl1X+TrtzZTeo+GmOAN9Tl+GcJefdLUjAp4U/VT4PnwjER9iU5hC2uzhbJ7ss
oI+J3TL9BL+AAy0TTR5sc8iD0G8Wn/sKTo5h2cnXqeo/I/j1VD6OoXDSYVX7xthkLrkxEGA1T4qP
6QEApUqzPQQ1SZUJEyQYDtM++3YOE/3P/QzVX3cs+wm5YOz1Vmqi8e9cLDJZwlv2CpGkkyGRU0fO
TOHVJZciHFjVJmQG95zRC8Mx8jzkGIoQ6IfdKjSx7OZGdOMXjUe4rVcFN29pIHKIQb+vp8M9W1W9
dPy5NIAbl3FGuxLLLcWXeTZqToek1opmOQMx50v/euJjtWKszfCpMumYcI20AmzxBTQzLeGDUvZk
DRXmO5mQsV8IO5OHHxgLtTcfVZ3jJ44vB97ny6SPDzhagBgZs2Vuj6Hxee4vOoZHkwh1Ff0Kjc8P
FatVFAQwC2lEW8a2zjig1tqIo+Z3BkT6tYIlvD4UHcft/M43LDf8E5Sd2dR1t0bec4xpvgWa1/rO
Txua3j2m2g2sVZh1lM7/bhY7h2Fs6BRhOzWU/4vPtYlqhZNbzjHElGG/M5lxzXd+OFPNz/6lQ1fd
0z97X2pUuQ4Wct9MJpn3Lx6paWSD9lFidv/wLx726DbXNEzVHeQk8D50FWvAgbF9P5U7zDQhW9CI
kPwqu673GabmfjlcUMVbeh1ATVuRLQk3WbK+XdwXbu8D1g9J/kEy0yH8Ak+1f4lTPl0Qnstu6L/f
gAx7168+hpqnBZ1oFRMvDiCzq5RQeyj0qYdBHWE8wNT9XIGUmSCRn2uOOAc110RlwOMJXrFdHyjz
EEvS2qzPE2D4jvEms6QRZHsm3H2Egtdk0VjXdeBrNz9ZE3YxJPWhHzxVxce7nqCFBgYh0hoyqdbC
DifovsexkoOYbw9KQfBgiC5c06ih3RLPm8G4IfhyawY49D3bFKjlFYbt7nQiQqqyFJzCcHj1avAE
myDYnB7p6/4ZXZ/JvTDh+aeHGiZtIHFqnRZRktgFrI2h0itdKnSYYG6N48fMs/hz5HjnbiZdzMYd
aSWmhef5ISCR4nf7mDe93LTpHFMMboAWRoXlauODSK9PEvkZxvRpBeK+lO0u48c7qzrm7yu1zVSp
/OF6nDyZkz4M1RHd7vfYvjEgow/ksMmas5qmYF9GXN7pXQzDIgsZVqMy8SFg1JKZfDX182Ljw327
L0nCm6EydAvn7MGBz1wu8sOAGGGbca51rcXTQQea0TvBikmzzcGKlJAZxhbbXB5Mds/FQnoQtBoy
sKmPe1c67E92xaO8Lsk0Ytf1ZrzzJ7CXm8zjTkNV0UIq/0IhDZJ7+Kd+AlDc0Egag4fNFGD1x6/B
M82XpEIQ7g+j0s6SIiMX3XnTfhfK8QXiFIkRu4drVU/3dDTkfnyw4rp2tfAzwtpWENxSMg6M+BqW
0L52cPYbo4rVtTMHaV48YfqwZSuUr2bQ9ZCzWcv6Q4MXDqyVrN/2rqDvXx2CwfQxFpXaywn236rr
jaFoNDPAD3dW2q9InPBf0HNF49HG6XlGbkQHdwyrV0TDkB9dDbI77BQDgILXBLwaandgT8NjnK7W
PYfYfVlLDt2OHr4SGOa8ibYwkykbbP8BcIwpmIKLulslMUuu/APrNPxRopjFjJnfCmD15bPI77bU
RW0NteXSZSrRruf0IVNUMajP1hG7EAW4bJcWKF2zbN6Lj1CUUJFOsdV5Ze8sL5ErSPiJju82YZDz
8TWLFiX2O6XDrRid0PrO1t49VBbYPjP2v13LoEcECXWgzYBWIY8wA5kl4nuM/ueFv1dWuESbsh80
i+D3P3Dhs3/ZZ4T+VMX4moxN8u5yJo89PxGr+8zVU8eGY1vf4ta+/L/10b4kilZeMWB+087luXt+
s3uveuNZzUDHp+XnwtHSFgf7DqjeH/Md0k6Zj6Rfk4QY/nhTpUaWFV7hmkrNr6tabrn/k8Mto9Co
YqhLLf9Www2g8vj8YG2Kf728UZ+sE6q7p7j/6AvuDzrPxZmlLdzOIqcOSt4Gk3yFzx9sGFnyQNnd
FKIddbDgEQlb3WcF04M/zzrr4puyFAYwVopnBKDx53ndITkqyRp6dWAEuZ4QI4EW5bdMoYNpj4pc
aJIblrLNl+2UqWaoQR4GNY/FufmuOpl3Vm6UbAVtyschuFhdMrwdu8gnUq8/YDy+3FKfkl13f2Lr
hTENpl40DjaKr6512zdEdIoIAQQniMu18bIlXfX55loAsr8aADolBEmJEQEwUfmNcMSGomnV3YkR
ajvFbqYYCN4WjG3X+kNNqsOgt1vmV49RcE1xTP69VyG/0IfiqOO36X8lydyaYmQcI0SBfoxgnBdV
iuM1Pph7LpJVvsqcVcGRNKoxFALT3t6+Zk000MyUlU3byys3jhM4VKkHH969JquBjjVc5CL5p1HA
lsWRJ3exmsaQE5TZmdYCASf8iizQimbMsZLWl/3dv1KV8AOfTac5ZhHZWa4zJbzq2ZOE5OX9TYMw
4kDv7tdfJzmA3/MWmz2Ee5PQdW85jwbz0pIAOPWnRnrTuI430imgM/gScLSHvDLU6w56QWiA/klm
WpywzQXPjNifiDQZbRfpobjzoBfCwvhCeLQSKz226HapZRpHzK9IchqddPBf5d+AI7Mvk6NErRpt
8pMDDyak8Q1NvxBxBaZCLna7o0aoCSy6CkJ4vxX+ulEj29o8Fc3FQ7R3EGTpK4FTiwyVEBLdN6IR
vZPZmbuwbzRd4mPUILjGTcJMeYAGlwJtwACjqkh1V21cPOsCSJM6Xge/huyHAtv3pB0hqrEcN/Df
OXYKwc/ZufrqU1bG2nGdYNgJmJ4P/WBu7Jfv4IVnsrhiUnfsunmHty5phBSBmRL55ZZmRW/zXbnS
P8i9vwjIuK8IEtT8CG0kA0pWfjH13RfQ2xW/hclqxC/C5PzFPC3p+2Wh+HBZey+xwprMtYjh2Qgf
55tBkQe0vhR5nPozRnSV5QJ0hJJF92s4isLnDRHgWdOvUo6/dNyP2TBmskRB4ywAAtACI7LJTa0A
B+I6K2hXh2z3ValUJffpzOaWOebjxXAlkenQMICHYM0+C7dQg8v52F92DW3JB+ZLLd2OhIdD5MrH
Uqeu19zpMgnKgGPOpysEZL4MMR3eCoghwzeR4kIn0g5lark5SBaE+F9K1vRMW0SHCMRpu5svaB1c
9ekclxrRUVtGACKe1hiQD5/HviPOFoUKZq+yEl3dsTNvvLgUkBsSIYTg+zMNTAQ1l9Q1h7a7JSvG
KMVEmHyAC6fl0kgbYc1rGpWOFu2ER4GHcisDMsCDIf3Ii55laaS5ypmdQ6h9EPBnaUbCFZSPNjnL
v4p38VHellQzd7G3vi66UYiC3/QzPnMfrL2jzIImsKsiiYhP7gWGalOrvSkJNgqy2nVvcF8Wj0OB
FZwU/4bBwqxKDWTZ3MnWy4c208hAie1wVhCbMFp/L4xNKc8L3aLYvWNkXNmxLp4lrVuJccCcr4RO
m7nXnR7ejz9vlmYDX7n0YPSZnSo/mnrivopei1kAZMAOHm4auoRY1Px3GYtMwVKGLrFO0FY9nJzl
uqNAbbRPQsCeIIn+fTImDz9BamgrHfubaOQpafIW5/2neZrGCnIY49znuz5lA2Rr8HvNNhVMtwYU
WUoqIJb1HVzEYoSzIE5+UM7iaoAnVlNrUjubUP9LRhntQgnl1GavwqWNUfxWgl7VDLLnrHsqM7gr
hqMUIoRQNCEgGrS8drKjguoBJyzsyrfUFre02407WTVk+b3Mok2JmEIK4btOlSM4mVN2kugeHStY
iXq86cpsENmufgjhjTcWlb85m6p+dGyPhrMYL6Nj736MVICAm9OK1/V3auKHh9002rISNhjC3yYk
IivX6O3p80/jn/GTs+oAv9056qMUZSoDZYgGlW3nAlqPXMgljMz1ZJnNw6JSoeAsIR8gFuBv643T
BBmY5up82yiSoz7N302CzB/5Q6hBk5ZIqjwwxmpPTB+sO4uVtzGBA/hpi+9FWNVfTZZyfa0Zf41W
GBnqSuDONxBKlKXng0oAuRfEusMLS1UTANU3IXHsbW3jL5dZRNFUccNHdK9VMjX1Ov3yS8HpNZ+I
TMKnMvZE7AT3NJQfVn5u+HkTB8XwEDBSL71KO5ZU9bJ/6GmflMSvCt1/nbMHIYhgzzIlEEwiNhC5
QjnxzDHg3HFmZzAUCavAHNKuhEbsYp7tnqOfreJSu9Ni3A4RnJSZ6PIHyflVHIeeJ/4zXSp6Qdlb
d80aL98abkNqs6gAqsOQ99OWEjncIaZunufcOKt6jq7k8tgh2Npev0L7TgaATsawZw7mGmn2dOlu
BYBlTEk8J13QvfLV+oHIAkQWVZndFTAjMV/09/Qx7PKTNRMlHsRLCzFzuFm0mSIP7s95nEVIJ/KQ
gcIn49z8tAyOw3HA2k9yZii2lfi9AJPlm1u/JzuuzHsjq6J+zoPXneIWszuhxJAhftyhVVyq6qcI
0RxS7lbq6xHXfWGFQuYyLaU4Zz5c+b1/6rFAke1MybPnJ8Ah7LE7+wmLbYHh07EpNoltoJ7zCz6C
bNdPZbzwfNBEeTiPnW9+2eIaWi5SQ8dOd2j7XbvwZEm3gObkARVe35D+pmnAy8btzpON7JqK+mCP
mb0HGTRUUS15NJ/wvaY6fKNg8q+LFzkgukhXZ6av2yAOKD8WabvYuuJ22VVN88e3rdjc4VmtnU5r
Ksv2nnky4sj3T7rRm+9TjInsjgx7hkfwdKrEcewXVpaDyHiKcrEKP9/J9++pdnTgP9y7wgE/iGmf
5U12qp7LW2myKpJqrkYABN47dIA4kWJ4wiHULyA783uHX9D5gHoFWSAKLV68Ih5TrxRWxVjCuC/3
7FEU7aPq/A22uf8jMMPUwcHxONvppt4jukT6x4tiuwRvfrmxWt///Vh1WXwG9XqG4Hrei75wKzje
YXebsth0SId8MISLGmCYba3GS0Kz46ribNE/FFSXJ2R8JzEy8v/ogNLmtly55IN2OrUhEV30lW21
ik5q3vLUQUU0Hz9wDsorwoqLmBqq0nufEUZNBuLLezUyscIdt+I4xJdA2MOY/KC3wQsY18T3c9di
/yxLNKgr9YwSb7Ale4bTARJVRRMTwDtluoFRnF2iVynU+XJk3Rxuna9MrXGGoJzp8knbZ3HsTOq+
80x3i2et3iQNWdTkdOdPZ4OUgYZFnhnV+4KmzLeISDqEZrYL78nRhmAdIeDCVYN4SYNUnxf0TWa2
7cUyhGq5DfCS9atxS/fKwlrXrGGhubq/2ZjOw36K1gaGuqeU40krAwgY0ZbvLVrKm2GoX1qKScjW
QgInfCoqZqWg1xmi+NBtDtbfOz2qG8l3QoWWAhEjz1nfbKxiHEedluGzct9r5jsl05qs0ccBs73F
P8lfXz7VHMu/T0ROcYU0oM/LC5t7DRdaXg9Af2nNyc0ELcYKiQa5cyexmqgTqkkGYgGDX1vKTcem
jzvZvXgMo/tSC2zUVFJHRfO5MJhCUVJhEJ2krOtqvhzuOYC9S+9mf/DKt6Vz+jcaBsdGHVfT9oKZ
OVKRSRxuNqNHIHuxNtmPxwrh7Jo+Cse/GB3H0Nz8+FLuQCuq2NdTw8V7ynJfnQ48tI2w6F8ST/MN
kfAd+/o+aOIhZU++SKqnxH599/H/TrcTpkZMQ3CoCzPPzSLFKs27U68XMFiRZopzYFQEeRTmAnNC
bE3ve+OAfCEwNAJbMKWimdwommkKxA4xdmpyoIyAs2RQy20f9YpPYjjYy9gKjB2Sgo0BtNK0rXLu
zqy40vXD66pyqjR/YwSHPyaim7fskyH7JbcFeqheRRw+dLceQmJ/cyhcxXGn4BQJggxOPt2i+xta
akxUdVjhnv6rLoNHFNBDzIGW/eimYN+YLiFmvu3vLzjutKMOSJDpsq5vJM3bMdnH6p3lG0XALL/h
h5uGdPBRIk+VUEXN6/ChMJMaF3byV5T01PqrvWBpQ7SFHLQC29PizbRQAuQuUqOnE8PLF64/IFxL
jhKaXHMNlK4GLZkBfUftjhZQdPq98LVszF3aUcEGGd3XrXhPtSZJHEac0TpB4n3SfIkHszGH028j
UKxyX3P/CDK4JSQQnN8Ksb97MXUG6YlIypPcdDzsdgSHAag2JWpdPpU1jf0SRfyPhDdQH49fnO+f
3p45i59d88Lme9HUtuNBNkHln5erY2GRFKlZgPmFA/5wphBhvLkgmge4vnegeO3+ddyyDjfe5yKj
oXTxCq2K8BT/iQa7rYReu6QlJVICYadXOwDPuYH7upF+j2MM831OWq9ocuIJ2hkkMCdz+3KL8mCn
tg0zNdtybLoHK5egh0lSwZ5xEdxpcDltBakkjGNeT2/ZW4Gum7uiC2gStMFv1Oc+HH3HbA8ogJG2
iO7FlFTZeWHZhYoFpnJTVNfDryCi7vR/cV2g2k35QtRyZssGvHGk4+3x4FGv/gRILYdNxxxBZyQ0
lczm411JxKVJ7qgnRfqC8/7JrbDJk5hebjMXFOrvmCkvJbvmLzTdqq4LJLQ7qsMN5uwfAGNr5u8p
YGn8PYN6SqUBBzCoTR8rxcv62Qy0j5JpEsx5exi5pva9DrLeLc9axvH/ks2v/AgZG4Z16rT9EJ4V
9tt1bLUu5QslWCPV0iL3d440/JwKwkHDZ5Fwhi3VWqmzIDH+9q1vCDQlZ5tZosVdD3nQ47kwxAJb
He6c12BgR3BfbTTimsDh4qpsHyXYwczJ+IlbPCKXAmYZRYSVSLCnzhfwuXtoO3vk/SiOvjBQqihR
S5OIOnht/gI7HgaYd705bOUDq0FmQreawIF+xYtRBL2Rxng8Gb08XNjZOwDkP+fqcZxCh5iv8vIZ
xF0VYCRX7ccs61e4GW9H+ZJTL/qUOH7jVWQYc65NGlJXjj4GTL/9bvVpME6OhWsJKTwnp03b7YH/
vCbULeqd/qo2JURD8Xq3PIwESWi4GkNqQ9CtZtwj84367TyhoUfpu2HMEmwFfq8oQcqntsf6WKFx
bfvGc5NjCETr/tyC/qq8qWJykIuQhj3cfISpVzWB+pS4xSAceHMcFJP5o7naSgxnIWOFt764WgD1
wn3KZHr6vci7KmnPt2pVk8DxfBMm9TfBfY3Tw4hZaB/90KDsSPQvd2yytR+jjZ4ea6+9xrQ/vx76
zIoA/csX9oCfCFhZ17zNJzqIJS01fN/Q+V1gRIy4E1O3K9+kA+3I1OFsA1C37xvr4eobhvWJCBmU
wngpgBSOtwAGs0rnpw3GSP/+Ns8rTNVwctEqDLoTVtFR9kJbtu8zji7UOTFVKDPouwOSpOrFxbq1
4a7ZOHVxPpB4ecHkMoStGpN7GA8VW0MrjPMbCdUjQtxRLPyJJJaYJB/Js34LXsnzYkGVKw3B+0ie
25bermbs3+DumEq0jPcJlTQU2/LWEjU/FHRmOxMhynphfCj5xQ7uJ/NQ76AZEcCBY249Jd5zSTjk
GssNzQeFq0naGqfcSCiasoinMqkSSbH32cl0HbH9ssmfP/x8y3BijwIia7b6/6RX8sfRcXWWyr+4
4fN/QLaB9MGUkmn2dzH1wD7SmB6xBOhDo/fdKJKxpY0ptZCtdMYKw8RICH4Bbsu6z3UxhM54C8l7
04992liLXQqBvbTgyvvPbznIBxpXmgm4JjSA5cRMnQ3hzRgjtfCjLkQvw++ll8LtmVz2JW8O5n06
MDbcZ63ar2FKsp6A6rPoqR6gO8u1/+O/ymdKsVuR0nfjzjZFf0egYNjIjrw/XZfsATqGgcNrJtX9
b2JFGKNWOEBCbrXCX+pkShYsczBwE0oCcmTfCBn0SoBpQiWtNMY/M5alCa9R00Kr8bGOOfIWNfWF
U0sAicLrHgTN8EPSbjnsanWeWQdrpgb1qgh3mCDqWPKgsHuQaEIAJ0MnDn65dBA0jD7ajdr/IE4z
b6nMXCYOt001TBnoN7qx/FFgk+4DhMmjbk5gQ2h0atNNhTkWIe8NN4XAR7WeeYw3iGNOptlHb0X4
AhVJO1bxlm6fVRCoPjzYS1jE3pKLvFM0Cq8TD9JdOZrJ41OigUFSQ1a4mYuwZRGjEYWFjrzLMppG
QWD8Oq8uCFELy4SsnIMXUriz2swF5gpxSnCRA8ett7sq47zhgyD5lr2X0RRpSDxZGZy5wrXSO4dZ
NyvPs2eThUaF0d9SsaTGlGxxi/ntG40mpLHYG0lZ2jUj7Bkr/vSqUZAnXTzFusf1SyyCHpqUYCyB
3HHw5o2LKipKxawWYPwAX1UTYrk/EVMiQD3PcdovHNrSezmHnald0Pbiu/0b4N5bbCg4Q20VHoc1
GMixLvR+jloV2P4GYnge7L3MkSaMJTy/S5hGJPd/74HTbJu2lWxNcpk8LmHWs/zHBokx5tAjFwkK
sdzbfaOk2QgsK491RLtSb03Lx21pXL8udY5jbuY+TRF8Bebo/7Rer2c/VgowbHRexioAtV2Xy4K3
/JftgAi9bQWJWxM4+aGy6wnOQcT66GFA1IJP6wIc9ONy5OZfy17g/EyBhCxRb+e4+0HvGvqnuDZg
rl9lbCM6KSp/VDH0N09oon4a6TpOLeN9o83vCYvIN93hI/WjsnO00iXpPAeqHh4DX7dtD43Af714
8x4JRrn2Bex2whYKX+JBYwBpiGiMxRcV8YAHLG2T+z3lukMJz7QISHiOROs3ZgpcpPJCqoYciRDW
GTKntqY6ta23qni4WT0K/DxszECJJotWbHUs21egJ5mqAoubBVpZXsTo+0JmZmrGrVDqNcRaNSTj
p9cg+NKl3WMk4KXq+ohghJY+/z+e5FKu5HoJF3ItR+0Wh1imVDuEV3kv9Jc/xoRD5Z84gwRgXiAJ
IWaY4ZnnSyjhxqq4psd6+jgt2VwNF9UphwYXKN5JBRtC41Aj75suSPLU6IjzoXDC+N6uX8DRwdnO
icOa20aXcd0Nl4SKLd6r1BNGu/QiuKepPlNz2wLSmyBo7RpkQf5TWCD/r87l6rlfIsZJ9l+wTX0o
ItdelFQLtpHS37hZ4/vzQIErTESMmhGLT3DzNi3v/y+G0RfbugzLStnEuO+EANP8EtBNMQbAjsmx
haPcqafLZp5xlX15AHio5AhqbBlU6U5a3EsYdw8Sid3xwQW18SptkshWglgdpYh3QXYnea8W8gXp
7iWbSNk2e+T6vKET5IJX/i4eR2KevlYXHpTr7BajkibdZalesobfW+Eoh4bqnaKJK1qt8I6wa2I1
mL7O16EAtjCMRazDpqK2QfOEiAWR2a9dsY7AQbcblg1/riGFBd5la6DozRzUmgo9H/sOfR+Foddw
8OS8i27ojVw6TVqQaG6z0gqrzW/eq6GmE/dCT7rWP3OtXIZmMOsQNDi81lezsqPsJiL9DviY1juV
3GfFPrgsFRWr2wWEJB2oQtZRiDs67vLzKBveVIjwUwV7CyB0hc0ah4u/lHfjb2A9z/Ov1+NI5B2g
oTWFfDKcCO0jwSrkZ5xIgY0EO8mb1Rm/zlLiOwcWaKpHqEk2Fl/9WH9Nl3SEAQvK/ZCau5wnCzAb
kUUIrcdZs60WCz32rIA/AXgnU9cFxFV9xngvOxmCWSzXveqQFnQqzz8K1oVchCB6+nkreolbiEFD
dpBhTI5J55OGPzVNl0FQSTGaVj6ctaknh62ptsM5GDrCBBhzDFUVYnc0siEreFkREabXcyTjlKXp
deeoiup1ovefO53eulryMISgd8WD3BhWhApm92R7OcS12CscTYrW8029J+leqBYhzR+asBX9lFN+
YseJhINpHT04t6U60aL1yZAMNtRmsi7ewqHIByhc8lh0lVPvzj3StkzEnJ2yOkVqEIs6VSSgjTfi
DTkOfpT4tUNXmJaI7dz6TYqtknt72fwU3klEP3XLg3srBrpKAUA0assu6w0E5bzQh/TsUw7T6E1R
FgyaGXgUmEeOEVOiQrO8IFDeey31Bv8j93m9siyZFBqfu+w2t49wQQjL/ZVkZF9zFpH4xwahc4cQ
hBiDd/ST2bM/oYoBMxVsmcUo2VRfbnC0DiZ+r40KK1qEov2jdsPn7mCkPTCzWmZrIIFb+ArVZx91
uf5jaa51wNV3NWmulBKNaErLhzHnTXFV3+wfzZlFwaKgnzerLiKvqdybPQrtOeKFsqrjEosQdVAB
a47wKB0J69/f02uigDssOiMXk7H+Vd0FXUS7rzX5MyanHslxdV+j2gaFk6uIsaC7YGjYDIiSYM0P
0+Dr+AOXjjjvdADAV+MNMtYmGiksD9nZTCiehjOBDfS5TUbI+Jzyb78vDer3L8H4S3UVIWMtY3Kf
JX3O9si0l86ergDQ+QvjR9YwMz0VQyf4lQyBeCkxPNWhgTch5x+dS6/lp9S+4uMKaqiJVcEuLiQa
PjllLht9vIatS4D/X0WnTvZfK6aNWGvKMlh81iBE8Sb5n6yhd6I4OJV5bompzksPxZ2zJxuBFtCQ
RoXLIHIxgdtVuM7dFN4WkJhMRHh13MQ0lCESFT1nlWcrkU0VqTF5cJeutwQpjIMEZnHTrNlRPnDp
g8+WaqyfHpgTY4OpXzGI/QgoORIG4SkIMV3ZKSh8p7WzHowdkvrfxEc+GJo57VhG3wjIPm+/ZhHO
NBXhf3b7ZRqtSY4a+9eDirI5bTaaZnkeWdfrr8NJYcvGOISoKoCL0RRwdZQVvM0UivPfUKDyY2Vs
Asstd+9aH9q7xHZm72m5tz7+MqNAeuHtwq16Kmf5zsApoXNBV3m1/ApIMyswpcSiH7cI04BdIJoR
ssP1ZuWgST4lvRScLjpj0iQElzwsEoaxn1oFq7tLrL8b8GSovRiaa4nHT7rdN+t+7fxQfGEtjtpn
Dl4V0xGewpmpBbUdd4G34i2dc8ohp/fvF/JPfDsCLOKwH5QV45aF1HVmhGpA5CUtLj+ZJ5Ef1oTp
nG2CfTcweFDruRLAioVkmkLgVuCLjBOl4QO2A6zpUPY5+uX3Xag/hoInHNkOaoU/AMh+mSmZjjC0
gElAuITEQofZLRhYh8cnYOMUVdKHfaEaV3EK702x0WnEtMGUKP0OhlOT3YbcIrzltC4b+zfHOpkX
FC0rfsGWJFpvhQ+uzS5pNL+4mAJ9GVXmKgJq5Rn0IXGy5C8brT0FAGs92FK4HIA0AE+ph9O8x562
NFkgIUh8J8YUKkND3Jp5Of3Sm4SsL/bwioGxxBtg06ur+bSWlWEMUQ4vlsek6/91eiMmvM2uIksr
ZYouJKJsogMoxv8RWQJYJc9CFcBM+mE9n0ZGcV2HakCBse8jLRVMsq5TL9gA+9anTJ/M8XDAk//o
qFDhOEN40QuNMcU6iH9EuvOj04QiwnaVnatgubqfkCba6JQ1SH1GuOYnDQ+4lw8tO5NWGC5XZmfm
OJIpj17j3GgNUb54KRM4YG78byVvlbzCtkjALD5IY3rLuCnwvc5iZpuG8NOvZf/xKxDHjuxxCMVc
W3MOlaI3mIWGh9K6jlDiRi2E+xTvQXbR8/IH6OD5XsxB8USrsjnzPZTOL9KIM2agvBbO/Z5TmT4V
A+J3tsUAlkUnt1lpadhdEGKl1dK7h2mQKvXG5TZpUwryXeZ6TufYfAmtSgltPFfT8rEC43ZiHzl/
DpwyE9CZ6r6C+75arnEQ0T+tqZmVlIiUbawjYeSVG9GAZQMzUDDfkTfXLgGTB5RLxuyLJjMnKWDB
uCjOn+2u5iIoig6Kya5RAg0KN0V/KOCL1jAzGIvhPbXVCJZPAIoJtQVmXIBTmMgnf9udtD+zkJMM
vzL+7aa9NG+MW0jd40ZW8XCyF9MldSjMIfVtUwm1bMy0zpg5H2wJDSIRfTzrCg0e5SHvk2lWwun9
RS8WlZrTpaZF7rHhZjKkrkBZVj0PM4OsqUc1up3MKVNKZcng7KqksfMcQQnRdB8XMIWnlRxdDCyc
pQf+DQY8ZvR9TL98ZTMNTDkLLrdzxSNZYU6jq4t5oxyWFYgyZ+IGJIvdClmW++XaIsXz1pzlZLmW
DdGffA5gq+aHit/1tdHOlcE4S+U9S0wwrsr23mHRpVNP5qVaII+zbQnE6JJseNhfZsidtlLt/b9j
NS40iiywSkRNA8+AVn/VlWr4HgBgTGIoNzBWFKfZClAT/bWZbBGD9f1XBv+oDHtLjJdE8z9ABbbl
BYE83vzkJGMn7OzJnDmrZs13pBEtFER+HDH2OrtxymdVZq8wNPkHVBDxIfjr8TFDMDmKmU/QFlGu
Bwxi3U4bW+tnsSpilJUh1eWJ8GZ6e+nOrUsOO0rNO1fXt/LK/b3Juq1JFRhgLHXjA82qzd7o3U7T
fIhSRdtv2b061zAXrPYUSmJm1HvLp1qmJegEuX02yZ5fdEi46ChRxVNyIcr39GE8T0zF1+jMQA8x
UrlkMnri2znQw8f7i3sQQ3q/OhHrLgoadyyjtFn3kEbhoEaErakvHKmIfuE+BV24x3EB9b0NLLJ8
S/B0i+qszo+p3QZL24FKcDS8nz1wXxmJNrc3zLGhfahUhP2pKxB+wbtRARAaf94HH5GobnNln+3h
fL30yL8inWGgDcs8/bzhRQH6rLUOcbUxfEuvfjtydj/wswNJ7OVhjRfsvr2/EcwhfJLszcQSU4DK
TQyJB43K6J/jwpe70NYPyWcDMELuQm8asDZHY5+BnkHPJe1XDxyNyorjdBYIUmnaDKM92kOVtPXc
1ffZXi46d36a8SuM/M9gkexGuwZrm7bCLNJWCmAZKT00EyCqrkc/6c0b3xoeB0YZUQl5/6Hlimi/
BaNkZQfY+dfS71gUiCDMFgIpZSsJoVIpJHLEz4DGbzzdWjPm6Fw5Yd+INyAnpFK212jYkDiASANG
1VPUWbjGX8u4CyY89/CM5sMlHw1ZpoyLwZTAn2ufSbuZwqPxlire2M83tM5gWrWyja+5Oc9Uik2h
WhoH/+LFtj184oc8i6dh6GS3Uz0XIoCpzw9gsl8Tp7T2E9pkjB2tr2y+0tls7A+SQp4hqFJndn9W
BZdUdtoojb//1dmIvpASSWxaYZQuVEF/li+Mm32Lj0qXG8PwB/WyLEIjA/uTFG4jtZOTmnu3Ib81
McimO368OimBwQzpRxFPfLqdFTHNWlmhMD7GR0FKubliY69wG+TIhAt6+tXgtIgu1o6CtFlZ4PQw
c4BqFqPdqtqBhPFaOjtSrQC7xnDHN+QW4EEBetjZEzNHpAM6V1ZGHvfMH4Z6qlpg3YQRPwOu0H+t
El2356R9jbqR4xh7XnOvlS9y41J/dijQ2SaGF1CD3PUxmJHjS+xOQeBnXdF3HH7X7vpavA3m5HjE
kAN/8rH5na9hkOJR49+1XjEC0k7xVyxUNtkpRDws6fR+yrpU9exs/k+xvaZ9ELXffClMITJG86qr
4AdMeo8sQcugx5z3h9dnHyvsxPyQ8TXcy4QuGxMEUlVjSLVGf+X1/JpvMR9bd6Aa9eslMyOR9AQu
E3LYVpdfepsOig/93hL86PhjJbT2ZU30U8V+tk2oH6HWJFzvz/NHNbYBlMIQHt3aYLabGVz78iYF
sX/u7d+xzF7xHJ04wpLfqo5zGunM/fvRwaIvSF8bi5vaG/sXm2GTQocvQKGzfTB4108jf+8cTmh/
b/Uzd4p4xnJ5hsPa1x4wDVXqFcXXkA3Ta7q/kbQxHJ/8QNNOLN636g+5jY7WGaBX2/TDIJVSVkuK
2GGuvSxRpvYy6J3GhUeET514mRqfxCGWY3/FgS5K3vO+cywih2x0BqSyI76Jb1dHuLpWldWQqmJP
Jg1Vran8aeOo9R4YD1lDzazQNT//mML1GPiodjmvSuRwBVU5pjulCfwEM+J1PtUlXxi1FqmcYBdL
kNsG/oQJKd/Ds9svh6SQT+n+UZ+sUyosy9YQnxbIiTI0Rsy9MiIFnIxLjUX+bo7pa+U37RloAhpN
zOfCzviQcjEDoUUQNIRAoJbwwFGSC85R4sxo2e7Sbhabkyif4Qh4NPkldcCZt8hpY/1zPAboiOxt
HL8rDOOP65wiYK7lLVuhbqKx44eWZF2FWKXLD8GVzoTDPqEM/Wh7nMSoaSCDAqa9ZjDKTTNdfWIh
8kbT2nmp1RZdXAfxRghzDypAgbIl1g8RbQNv4Ai8C61ykEIsgoEAIJJ8/YkfG0j/h1W+CPj1o9xx
wEUJEFkm2cvA+wf8bpwobq9AfyMajGQWZUbTfG1ixkb8LiUZg0FwoGfF+KM65V7Mzyi0GIQ1TE0G
ADmF2c7iWhNBVrSmFefzZuS0u12Qk3uxtBdaVRniNY5HG8HqaieUeF7ZyB4f6z7rHMzmUV1MhiYm
clj6OenX8E5UstGEFUkqxQokJ5Hx5LmPknMcp625FcQRF8gAAYa12Adho28y+mBAmVGU8XXpf1cb
xnARestIETN3CJ2v+iz96vECwON+oRBC/zVkMjgIykkJCnjAkW9JOM/zBFI+NJ/b/OgV1o7dgUZw
alVtmlkkm1MdX00w5cqSwtbDwZeMDHLCukkejFMC6JXCXOZc5pLvACxJWaqDPW8jtXjTwgo8ooYa
lRc7U+wz0QrUSsbjVBrvJa+TukY2eLwIwPVZdZBHyyO5hpVmsEWE5csAhjMpqKgbqE46em34AFiM
a7Q1RfPsYN8iCN3Hd4YdYc5N6N6eYJcMlegvC2huo93RswB4fu+mUwx+/L4lfeoJ+QXCLpZ6w9RR
g2AcNUKKoxlagpnTEkNA6SltZtm71nQdKs3leb44itJsqQ2/gNPKq6hHKSjKMVBOd8PlBeBg9Oun
aIeiBYWhNU/engdxs5QoaqIi1NlBbxTGRFCp7ljPVSVfz0PZpKXEJEnmyqUCzDd33vPByYozWZy6
7tYzJlw7Hr5wlE8l0PZgV+ZjMguRbQpTFMuBfiwFPOm9z1i5kZPUYujJP7dGQQKadIQuRkJDpsup
CRtUIYcbHimmNx+mYWJI2lGHs5yTicjrtJ+JA+wTwxWr1sGeNLXPUagXOECsi4bTTGnYfa6JGqoR
9eLf419qdQUgg73PoMAurFiTWqb0r4OlpzYWwu0+rEdahRP0r1CTFPVoadQi5KEFYQ6i3qOjOKAC
fCX+Y8u2G9XzNHjrhx2mFBvRnOp8afgB2mfg7DK9QQ3HefieC5hajANX9/0q5wLzcx8qSWsEnthf
RkQ5Vb8uW6+cqGsSMjaUEJ62EV0G/r1DszpbfjNiyBar4kKqjRiHq8cCmiP9CsIBTCT3QyZrzDsT
KNtK3Y5GagkPbBo+C/BSQ5mVgGVrEi+G0HoWWqeZwyXD77sNikkD3z6LHyWJMQUDOG5CiJ1dDpi/
H66Jikcf5eVO3RLl1ZGhf08UZKp6pNeeKOSB23K4ykgJHPtQiwfj22VnTki1vLfqiUyCYhIN3gdE
to5W2wL47wT1EJHitbg44DgYwymuMrInGT443oW5UEEw16IbR661M6rU5/LMo+RJVHxAFsDxYhtF
KYrn/y9V6qAw8FF5Hum8O3Gfl+k2oPmirbol2xsdXBRr+1lPo5LbQcM1twm6RkraFXueg/kZZ4jw
T44ZCQXKkEGs6fWBX3OHRmCWxAVNP2BxCjri1sxbZTMBSORrPWtqeMcQoPjaPuxpKOBvPwuB7T4M
Q2Gzmtvoj5ALaTn7RpUY94obuzRt/g8Fw6Pf2ArTbWnvQkbhNs89wwi7+vynmhr1NF5Jhw5RdOj/
p/eMIJ4aevlC11ZA6FKK1uki8rXn1db/JzK+EPx2XVvSLNUaUs1g3Kny7ea1LJkI77Yq2y3WCoUY
J8IQ5eE5hxac4SO+vZpFnKPN1a0+F0unvUUlGgSQejuL20sPTFQ5Y1lFaZbMjWAENd4FOSWnqa+m
8+BWYFHAXejXwRG7ag73W28LJS5n1kTO81CPw6mZwcaUCo/U0Z7HJs6h8CGkOFUo2g9a+ahpBVI5
NUqKcS9TuEPdubMvwgtQwXmHgepIe2DsY3Y9PHZNcydEoI/Cg5VA+hD8sYyZ67bTD2AtfcMwltpb
jSsn0nVF5JU+Lui+8ptMPYX2un6RQUFKKQPLyS8Lj33o53KfpppCboFx0HgM6vER35z/jqfpEKdB
1pIuAcVOifbZUAMfSIjb4rJ33n41Tb/LzV8Mja1ObAQfgqRS1NHuZzmalHoNwoO2uRdVV8rcLPJe
vT9bXhFkozpwwCguaTG05Nmqi6fZYQlv8Bg62N+/c1L0J5loReU6HcguofwMetqluD9tHJzZ1Cto
Gvi0/i0I+5GnTKzTlikOUb/if/KJbBtoHtOGMJvdzpafGavdMdjXOzReEAHno6yyoRk7vGLBChvf
vKY9wZWS7sRAVIBVit35Ua0fNFQarOBcyJa9OAW+RIHlFHoTVrt8ANUoPLL3lKNQs3Cw+Kou3YE5
KVY42RNg9sHthK7m72Fhlb7jf60SLXuHK14+VC3H3522qjeZNPSJ24SV8mZ+nzj5HUNKdyBEVVVq
4Y/xIrGAL9ZP5fi7/D9s7H0eS0Us+pD92pMGfAPxpfCmkEJHeIcc9b1qcaEkmQ31+gayefR+AeQS
fZewZ/WUEzL7oqFX0mS9x3cVNLX5rXWtNsKuM9Snmlq7AY/cd6hLeB13YnygxKLKta7/npyMAjC3
I8PC0QDxd0NHjZWKr+p3beGtc/XNImlPIaviW3CywNb+YznTTKIiM0qOagbBM4ItLxisSHPpJBFA
CtnpW0mRe5wZLkWuFV/sT6bf3YwXj/T/wP5av8MPWBnrAMwmMj5SoZRIaRRpWA0LS6t7XyaSZui+
luQnkNGQG0ZEaOAekaoyN/kTp2hi6uGK7tMHvVTD668kn5OQ95rdQMGYy4EaGZqcmEawiZrbqdQA
vnKBZhcV2B8bqvLT4YsjArHnzZeWe/ziVQfchMlCDmGpkEFvW3UpThr52lWvHPCLVRJBxM2PMkDF
1CM+SSUd4Kkd6S1WnHZyU7D0moducSMqfXxWWQT+82DsfFVC/bIKyCesu71X0tbe8nJclMHmuWfJ
Lx8zjYNeGZK911S7eURczIjEHnKRXGLRL+gSUJiJJSQJmXRnZ9SuBinEkDrle0a1ZLvZ4dnhXc8A
tkrnhmcP7QeaZoBOncRxOwyUqKkELpIsdm0fEQguef19hynsnSCowzJ7YMRare8MuA5PI51eGCKI
83ONuGGy+rC/6JGgP/SFIdeXMXkIWiVB/EcMCkySoTi3Ss1dJ17p5y4BTakLSxvL5Yxch0/Nnhqv
Djj/V9iot08kar1/7WUSiwS6MDHfyRjX3tkH/2j/r8LiwKI9XCMDsxQVjWBFea2jmNzwzhN0zN+d
wz0PTyZQnZ6dzvwEbPNf4YHEg47HkkkoT0ouKUF8ErphcD5y7lZusDTrkksfaEm4HZYDxHCEPas3
Dzllcn/E9daXtNAxHano337CfhWOysZ33/hZ5z+PIjsFEA48fsvHhLDNLV7nll+69fu4TyvA8Z6f
U8XceP79wakuvZPyb//S42oP/tcvM9mFS3yIl9yed1xGoqchMfQPyxjlqKEs4UAsVncdmIHQUHTy
HQfbOpF/MIRORV0a/K+UquacMU4GmCPEl6CTott1UnWVIIbH+MCk/v5u19FSrj5ahWu3q42yiBqa
TViYb6s1lbkp9s0px0TyNEZT0LdHed9Kara1FjwJflERGss5EBAhUP7TVizsmAd0+1X83P7ArgU+
x6mP532sV5UuTfzxMxUd5LCrRBeR7KE7ErnZGjldUF2R27fC53m+1av5f7ce1pKYuNgB8471utIl
XMNHZGXRoG8c+Bupovg0I8bwvAaO3/3ll9wHmF//DKf3fOX1WaNdl/tkpnbUu72I/r0PiWwsMuQy
KynDp0nlduPOsOvtSXi7jkF4JdV3wFa8gEIvy7RBk+M1tv4rlBjFwNQTw4H3wWKa0TkuexSo8VLr
NNk8UUNW8stbqzkdtguCKochf9A1fxjpDnfbT4x9C7TAOAxvthkAlyCFyjKEuql959pKIf1v00Hh
llX/qHp58TR10KdyuBwLz18GYhDEqqjWAkf19er5ReAHL6Ham1AStB9UAy9qqTMil01Oi6YCrwhS
ni+5QAB7kX+tcig6nNbqMYCjiYju0EDso1dfcXg0C+KryZG0s66rOZK54vu073iRnApLVwfQwMZK
N/V1JQ3V1xJYQ683qQczUdzlsxJI2UMB3UlvBHQgnVtRp44y3VhdkS0hgDEV3ApxjE7I3iEnfSoN
rGX0Q45W2ohMyBuTwEslebLE6n/5UFcuTwK6u1BZr7I5GjBUHsTMAlt2dxDRYqHbIM2D6phe1Quv
YyUpwnK89iFSY+RKu4NUcku4LbJ5z9RMLfoLZhc+R1FnAaTUA4+Pn4eNrrQF/DK+7P3CGN3CwLSk
3rHk+R+IUWvYGwLbL130gn4iEsFJkQpfq1uAz7muPID/GVY61kOvXucXlaPv8f8vLjCN/NrA/ICh
DFVRfyyvmor+oh+etk38BtcCKfIXE8dMThNFw8+wQJFDQEODqgiGyfgOJQC0h1tm0qY0rBjsoK3X
eBl9Uj5o/bOFGu7jinhwVUzwhlp/ASVa93aI9ELyV4BRedq6U7MP5weTT3dtz0gzjFXfDWxEu4Mi
9F6Lir30h+z+3vZyOaVrt4tAoPiHLBN8lyFlqgrQLF76pEj8lTgbQug4YPGnZVRujCkpY4Gcf0oc
8j9JmihEsJaU6xtiVtkF/dVGwQFhyMpJQ4xyd6epKiyOOGptgmEDRnHcejerHQdfIoR7m9itPdmH
T29bt/q19jmcqk+caWoSAcguenB6fuQGMHhKq63pVy28llAuNhojlIur/5F0X3Mw4ghuHfct5zeM
w5f3M4mEwigF2Th5KOJ3Miy/qO1cYeE+F/qJK3tO4hbk9ApP5iNmuinblLO32sEI77+69Z/3es7K
SK783sS4+xYQvmFO8ikyoHTEEdwTjXiCFnCmKIJdOa8Hc+gUFklMhb57pg2h1bXz7K3K2ptvU+hL
kiEubST0v1SpyaEFFQrss4b7QIHcUI2DKIAyyo/fh0EolFE98Cn86RttGhFq65K7jGQmsfdDwDpB
a6FDKWOXnUE2hXZkH91+fVTOV4bNaPQKXLzSzIn3Tddb97l8Wii9ZscD4GZxf/1Yoz84V+wXX2fJ
SkEwTcIHeefez3N/R9P/85B+DNm/WkzPoRhhL4//HDEeYaJyabmEhw5W9cR3p/W4sj5vSdY0vU1p
kuKfecPAUubp2togaewoaA+KldNipvgW84tmdUiE1bLTCsg03Y++xz5dbP5IJU2KrgGl4JAkkuik
GSwNso4LRDvauBe3MboI2TyKwVadzqU+BW0zzboQYzQNIjXbpFL7osN7kDbRtn3sGNUEZYhXriRz
b/L2pSITrYc1kJmeu+VpD00wsc0au/XGYFnF5ZgnIv++xcVUTXigakWDe7M/hKGG3CFaskZMJ/TU
0ynrTGhKf+Du7H+U3RlBpey4SjsEchFKWruoRrbODu9+EWztSEGbxOrx7jvY5q1RM8opzOv6R7CY
1APHD/kiSKONU0Yj81OBUlD3d++9k4M636Cg8XgDm8rKT2mBzgiBp/0PPyvetmQUAEUS5XK/QXEn
FX6TD0ESXZpMz7gu97v5V1hY3VgWPabLeaCBdvpLPRnV2952oQc9E7b7L9khXE4Muuw8G50/zuW1
z/eNFG6zGWtnZvW3nyFaAYs7nxJCBEttxpZ6LkRwhovkHwjixHCkchx9a8PKJwsGkzNY3lcFL7Kb
u1zskfjeQ/Nd3kv2fM0n2FLkuppGTudqi7EgsEBc77fdK8psLFUtqL5ZxlAk9l8TFHqF2SLlAWcA
bzwgyGDuKFN8vRfbkydFjE+DPhI6kVAi3PcG3jT94jjc5mkdLbi1cRqFehkPlS5+oDU8eaNygnjm
tXgenRal/sewQbGHuRLH9Tq91eMhV67K/rcYXJVUUtBkd9AClQTEBM35RMSfOII8hk/23zRAuU8+
W3TeD2dvijOap2K2vj0wb7yhF8tk+3pwJJn9TNALBCoCbRLJ9+pkXEqkBYmzNotCq8oh9J3plu0V
8qckW+HFqISoc4qDOpRc3EedyjmI73CPRg5lsev098/9nA2jiShrUBmKOXa1+/3PwzlBNs8JYpa3
c+A7dED5iYiTpgoLE1jjFkHIZ744GFzORuVR2HgAvwTuJLyopll/0arp+28JxXn+Y8TcWLqrQ48+
BS9zUohJz1d1BFlnq4X02gwvhEHqIPFoafary+xz+MfYaD/89/0Wq3PA/5tD8S8srKcRy853Wv3H
wv/8r85GawZpg4X+COgILSQLQKLS0D3gchVXR8jdXCfbwe2uIXp8pPmU0vombj/+q+EEIuyPSQQY
UhNxgSlY60UIAqRjYPcGJaXKXfOwsQeQG1RJzIxPNEBXBTK1zH+gh5MDT0IpFn2xIjrLhLftnK/v
SGzfq/oXv6ByzjgTzqvnNVXsZ5mgYmTUPDMhE3E013iUgu5dS/A7jrEpcmNywbBvZ2CaMSgDD9qD
KX6j5CWcHWBQVEvS/XnaCQkWELT0QDJYOzkVEtO6XxNDPqBe+/Pfez/CLqQHqmxHKFuZnzghbKHQ
o+EtTlB9c6xVKjnJ3dRhGZHtdkl2a4V89c5JsKipiQ1GMzPvzP9/UTfkXKIJmJL+ddAkm7wgkWhG
hOHdsbYQ4pB61VYmUhCkAnGYA4UKZbyslWDpLzMz2LQFEZ8NmUCtCcTN7GYlyNByO5wGmXHL9Wiw
I9Pl7Lccskp7DFWQ05L82Lk6B8LCRq4FirBZZYcDCUSDuDvsXrKa7puGFxsLTxKxwmbqgFlZqJU6
Rnu9+jGUyGdMhLFFeUG1Zoi4UyLl+2IsdHSWJ5FZh32hfs08Svn++JAQM9h4HbhOyJ02yMPtjjsT
pziaPCb+c0e9JOe69P41kuhtN/lFtntci3VCn+TG+mXPKiLrw1SzcK5vwPXOKZFcai7XNemTsXw/
78IGlOqphNNI9lVtCakjrMeGRoaOQD6ZXMOsuJ3BxUJpBWPIFilluupGSQkq6Q1krm39PI7EwJux
GP1OyoXu3TQHWeuwuzD59N1Gvk6iJqLvCKqyMo1UZ1bbM5UjslI3tA/C2AfTBVEFSlX29xauhjuK
TxfT6xW8h0+5jt8+g4OkFgtyn3Cqlv5lyKF6DqrHZRGOoBHPYqdzeVzBr5scJf5+iFvSt2wkOYL2
ODO+YQCRBRvnaHQ6uxMr1F+Pg0qdEQtKUiQ2PylDbjCYvySwLCjJfOoB3q1nZOXucJXdLeDKCmiL
BNHuXCNslNaZLln7Wb1Y8tUtUjlkjoU4gFk+5D1rQrYlyLozECuBaQPzzI+yDYbvRZ3JjIFNnvzN
xNI08zDIh+iTOIvSK/PTb3Pb1tVettMCGvFiu8yziiPXzmt+bbmBjlM37mZgf7QtfYhotOfuGhuy
1k/Sa4g8oylClPrA86t1HW+a2SvYyLaJK9M5n356NXgKsf/zhQ7nEn/HcJ/ZCwt+V0i9hZiF2soF
/rRUgrcaAm3jI6PvH73HYcYTyqoaySn1p5X1vqwcO5aIyQac5tGtf1HcxqOJCpO208f5g34LRwFb
a9CxJSna5IK4cMY7lEfpDbBCdYsp0YAyBnS1lDa1P2IFy2KUQdLiFA4H8iezRC4XvO8QSInMH+ax
O35d3yrRZEhP+mO/QUtmhuNOnY3EMkoL7ePqg7YiqNtNNY0fhGAD3iyvTJmUzOqZQtGAY9v3zmF9
V6xHtY7rx5Jsnc69WZ/v6+49Vz1XtMfr69ANYyszQT4RqLMmoSJydcwVPo0qIuvqzCPlmv/vDEH4
X+F4AsVBqhRzP5UqdpVGHIXmOA0PoyCeHPOFJ0so4MdXhb2Kq8usX/LHQq5JhskzQdN5IIQw60EV
3w0UAyLjqwTZV8K3CB2u0HbklBtDIxDWik4NOVW0y4omaOeIsZKjiBpQrMmAXEYBl6Jr/w4XheRR
kIk7Xcjcw0lSvwEc4Cnc5b591mRldOENf2ELTyMOOLnspc9UObiLrc0SEUlOen5241ns2WI+JBsH
c8xlNljXskRC4gMMMaO8lsNlCOg4TO+7oD+aFlA+AtASzP/C4FsEfyisuMJI7bz4WHMTJ+zY2UGz
jxKZFKkEkXiu54YoEMse0a60xuUasd6qN+LT4INrATMZpu/HStJe26rdpFgrQ+lsciRfrYbxK7So
yKY2RLnZe7jb4UAXOlbdWjNu8P+moEb8KQlSki+i0qRm0E/qOLi5eBL4WjaFLz5YPVy69D/VY/GV
rig7DIHkVgIK1TtEwJyTrdyU5d+p5FSj0Jzhfubzyg2rMJqVTU7kHlnR44Dsa9y5pxmzltRXxnCx
AOtRyizvbLlwn/eLQveHYTj7sWGaG+bh+ThHQWIjL8XAZwEq9XKFxDGFPekjkIj73m6Ye/T2keGJ
BYhNC1zx1QWcT1gp2z5In59hZ8gvjXm5rQVk4H6MVGyexCCnJTmHMJM8vpTnVjsQ8hvScnkm2Asb
/KFzdfmoEuUXL0pmXOdCAFMovlOVL41tYEs5kHXgqNkG6G1KpP6fWabvNEMx4yw8Rs6tgCOG6DiA
ro6+Ui42AGuySIapleUI57QN0fYV0vNVy5HHI6WB5UR06NYD31WygERFdw+3za59IJZmskJIXM6O
ySD61VKKceTVI2Pgod14OX0GZ4ONwXdNHYuEN2Zavyg3Asmz3JEVeFUENe2id6gekjkc2LxJp4Jv
dIYy90M3MvnNMyI+Djs3aDAcKi9yaPuTWuYhZzYTkv4TT5dFVTuIC2oNxWO22097+FGdnmFkOaLl
spbIFWfqr5Y9g4BZUXBBkn+Obkf0lPrZhfbyIO4HSsf9I0ov9inmyu3uR58L82mLOaFVJgokHQh3
/PjDo1Ssh/uUCkdC9LOkakYKv/3+0p8vRCtXZeHsC4pihp2tFr/bGFhCo/pR3UkNqkTBs8wl3GHm
Q5qyWpO3m7rUFNBUPqqHoAJbGvCZ+/cFE15gdKoYVjO6OJvUp+1RlLUbyFBL/LAi+z38RDhB8IyE
HdHNlpJRy46HJh5cOa8kbO/rYk8CoB8COdsd4JotjCzyL4Qc5NJhR9CMrZUbRETH7Cbd/fdZOSJd
PIUe0+xjlHHB/IRC044X1U1FBlEIEh6TpvbEx/4C7EmCFDQouP9VX4RqGHoEilDOUE4RUL6T3/T/
Eot3Skd8+yxap3k6uhep+ofrM58jBL5QM/dFhplhGcXIkkgwjR+nEI5F16P5GIMkkTcxt6E9691B
nGRXJafOlSrdc0zjqlQtss5J22/KTqMuR7S/p7/E2LH/2lQPzFN+Mm0L61/wWx8orQ1GL8oRLFmb
HzNod3qa83McRhrlR6w1W7WYeu95DCswbNVra3/V6TYqxwabw17QZNAJ6LraQioVdh0pgI/P/Vqd
+2XZhKANBJ7/PzELSM47VJv6vNjyGgYNExvp3/JE25OIKvHgRFtmrlbmWl75g7Vb5GkcrqtXh39B
PYTSiOxpUtFacvwvpu8sRvQMwqAaZ32JUk5DaBAgkRPY6CSNEcJMKqiyfI0iXTAQIhj406GDw3ds
VZFpno7B8DH0yiHcul+8IEfS2uoYHosLYmcg9P5KuwnT2Es+i+xJzm6qch9SNOMvoinPAxleQCeM
hH0+umBwEioTSJUlVE9oyMHIbalsk00X7jvnAMriAjzComNdihtqZa40r73B9enF6XPI3iRWDzEO
HoyyKgfoZ6kvPpd5JxZsQvZQf4rGwYBk4UfOEyeQWCWW6B6TvR9SO3RljO2hXd914ejn2PwBCGKr
sM2U6hgHmeVAo1S5TIqfopT5KH1iWRpHxucmswIdjlnO8gGUJPJHxH2+6XoPEKErq3Pi0GLdeU9w
E8RNFVB9GaYFqsJd1FZ/gaBzZDVqt7hHVsx54bTQsSFJ73q1ZuPiJ/EDvwYSuKkMAhaBFH9qTsP0
VX/tkhdu+DVHOrVCDkOha5RnFoFtshje9VYqPv7ICp+nlC80q0qM54cxotab5sQ2ZPWWXsB//VhN
nS8VNSF4TOOGQQBupTX3VW9QQW3hHDIHOUonQau2rNysHfkwhalQxRWpn7T3jHrQFnSHiPoHrsWh
uynbUhMGWWQRr2omaM25MPCng9nkk+gy4JWo2VkXzq5vZ49vk3fAoyiTvLgtUswp1M3j1YoGHJP9
WU+d4GdpgvZqy8OnFV7IQEQ2xqNEwCULleMFaukTdGK/KhS8pJN3etmeCnub4VAYkYMxGAyzC/DJ
Vls902ISM+/ZPFhFEYtyGa7DMYNEXRJLtXdAkLqLv+blkxpfDvFIuelFxa9WjdPrDT6xbf1ZBvQY
3nFgCAcYHEMFpzHAsea559vBpUmzMLO4Efy6lKRR03roph23aOBqqM3/ejCPvy2JMK9Tp1lZ2uD2
fzuZE5I97/KoEutLX9+Mda6igPRwP4OGP/qXvSMg6AHMAxzab88pN90jYcSibGatkogIU50dp0/1
QQwgm9fQAgaGrk9wIfBV7PZU1e/zxhD7TzB6CYC3YkhJ0VXKtdryfDKXfKyERGQS8hiYU5alM+Lg
GD0J5yTnFcD1fwL+UXx/2CUuBWLf4p4MdjTGdb+/iz9UzaaQQb7Cxa+SJ84BYsD9ewobbaKw4YpM
/KZXksDTN3o337g2QYSuK/sUDIycgPg7aP5xIMXY/hdMqJdIsRA084DdGfwh3M4amR5jz0RZUq60
7qo9f31gbOVpr0YwlFCyJaBq77IO74UyoskwXLRtziPtNKiQa5cGh8NwvVUxpIv2kZxdhRxcrEyR
8U5dtHtCFROdrDEl3WDv7L5MXWV59FfwdXJONCwcSsmsG1MHZBpSbtNMna1zPODG3XofUJ7uExBo
jcL1ZUZP/tPnvfZyKudq6/vZBIAz/bEyJDF3OEVY0+4KQOStkfP0utfJ1ZuZCT924ydFdzgfBChT
xjIZ8TnbnxjaSfLm4uOpAiBQ4RY998LfGMW2MCEaPrgxSyUrA64Mn8c5gGr3DpOO031EsNwB3ZVU
U+piKRwODk0+W620DCmM2b6CaxV9O0zB6yrOXeyE2moto306PrPaZMwszGwraTrwD7m0+sn7Kps6
I/xqKp8Ufo4AZF/OHTMPboEBFoJH8s+NWdueJUYJfmG59ZedHOw2uETRKiihCvtGnHwWo9HWF0pg
AdXbvZQ9EObPPHn23sXRJQS0y11Kfep0NA8aT2147FnMTC5gcOfAiGxowrg/ypwDegPxAumepEX+
QVIFtumVX9WwFWMBthgVsGtWTMOXXzrRT4obKcLbB6juCbfa2A+lC8mbPwwj3m0djMRGFzgtsDxI
1pjQS8CLmNp1ukpD1gUQ4WiQwdnDpQds1iIc64RR7H0TEdYRYS9fbCfQV13xPPUReTzVwCARLxwB
LOX/puWoSnnVV7A+uiWMRR7Umqovn9FokXqUeavZfh/IRIUGOU1bmbidXvOax1wzcvSGF6ehXpVb
5ZHPQQ1+sM9YYaDWtOkWagBxP+SxVvm2r3/tHbDiLyi23LwKzOoa6jH0ZTJ7tZxu/uqjL9urXwc3
NKztuTnEhxMiTUbKq/Yz9lPgj5ghrmhcKpU/ZGC71+HGANmB19mmmarLkwEsBsWjUi9ZpFB/Xp+x
GFn3q1vGDzFh0zbd6Ubgk/SnvluDD3KdT20Rhjso/Rbf9PZ0+pwG/0JEiOsFGUsfcPjFpu8iqHIy
d9Mz2BGoWhNe+INSVNW/I3dBSfS0ENVfDDj72e12V4Qs/N01zWsNQ4koDQqBf96xVAVxhIQO3yHj
XvDDVMjOnkiugujOrKOSBrGfP2nu3U5rnXg1kHUrmbDIrKzVHyYrUfDoYnZksHnislnjXViC7Dwt
GDdBu/XqFNQ6opcCUbJL0sdFFyYcT8Q5yMly6uu3Nl9/6dsakTBJCSbSTgRVN09fLpYDReqQs1Ur
iIaWyrqrr3dsW8u//8SRvO8mEo9/GQNg2cNvBllDPbLm3+Gr1L/QxB1hPEncH3VCdDHpT0Rv8Qtt
SRA4tWznb5CJMDaS7DJocgif6KP+jBtH1bDpaKLBTHTdq6ONl8KQBjC04ljZws1BJ4E0b6ReUDZj
hcyMpSNSU6EcUUGhcPpm2OCKR8LC8Ck0HHpXs3oY+6qgKiXMneTBtf+m3R7T0nWGq+SPebSByg8K
mMGAAYnMvYWgBrRshGRZ6XgTfwkL1Wr2diyd4Dsh05JyQ+QSr8lTT87tx4krKnCYdQwxV1vPI/wx
ToCdnKMcQHpsYDjsRE3jaIqLbZ+miZbekGhk7qAN5vzzcmLeHA5Ws++H/zx0uE7bIZKSL/fxBd9b
O6wBpLE10Hy+2++FZbPfDlkLZKYt9WsJ+NyqbQrRkgeKC12LqYuSO0orfvC/hIJWa3uXSMO/nyer
LDma0fPPrJM0M8pB6i91vsFBZNzx7PO7UYbptvGlaEnVin8S718p2DPbAagEza09re8OaomUTW3W
wI8M6DQb3a3ARH2u7MwJMCSoMJrMBQzVZVT6SpcGvdMna3lhRDkLzbhdlxbZgDTweLf0V7Iurae5
ltP6YbpSXXqrbAT3W+UFZSHuXqE3WNF21jEOPDhOvvHc3lCwgOH8yiKiGYkm6OooO5KUFytJF1St
Wh9OrAEZKlMnFba3e9AtVxU6z8+y0VYCiAyzT3CsdGRmvYLyJ36u7cPyfEpPdIcD1GRntH0d270s
k/Deygmi9wMzPXakVUgx8Vbb4ExUEWUYooDezZZiFIhtEWNt1Vw0Zhr0c4KaNvo1xQ6f2Bh+Gc2C
rppcYk7pBNYVuTMpf43bxSnynwW0Zy5/sx0rBz6n2JXtpjXG28xLtwrn0Dz33vlBV2P7sTmR9jxh
ytUOD3tdsF8M+lq9P/A6An5Une3zoqWyMnhVGswnWecaSmbJYWOJtkFoTL0nL6jNOLDpdQ4P7f0y
XDxl8KufTM6piUW2nXCflvYXhylSj4p95dS5F2ZBaXvtGE+AG6HrkoiJKd0hXr+CAYOeF3D1DCul
2s9Kvzb1hD1VZzEbzvgdAycbe83eKvSfzao9A2luV3TutZnxcktw/1swj2WMHP5a4TjbrIbPbZd1
OqJjVaYdAErb2N06I9DgrKCYhg58GbVB6BIKIkHtM+c/iDPIBbvOQTzpCZiUO4cy2AtHTUcZpT9r
6wYlv58SzVRrYv5btHLJWHXzokn+ZKBj1bWy3fd2vUV9YpfbTAdVD0MrxXrp8UF/2ahZ0s8YIWu6
NWJ+y3zYUvxN5eUdeMuK6V1cNtXKDlghjSro2o5C5pSbKuNsBXaplGCZmGWHEGnolGSr2DgrPT4C
OsHDjr6BNQZHqXKPMIxNZ/ynkH7ke3x79nT+kFJX7YzOUfLChKfZtL72sLVB2DBp6Xy1gMbCZaii
b5WRdQEONCtYxZa51EwRVTagPc4uhfvMuGED6C+4a4TL3lj+9EnQzK4mAHfZBvmWBvKU3on0kwRe
qkYLjh+kKMj7BstrKZgq69ckooq+RL5Y3moSR3P2dDkQ1Si7ouJuB6KjRVa4iX5sZ6DTUl+A6e+f
uXVy8tCrz4dT8Si0xe3QzCMn6jDMsY+vyNodttyaxGHNG1F6puP6Q8djNsarxXLiUxGRn2ILQ6zk
ClU+1WQclnetM5GNvI8AVYxQNw76Nsr7Fay3Hm/mmlXmNKwVBSYWVOI0rzXOHJXZ9m31CgDWnuCz
2FnSHhFDEP9yoeHuveCjw2edYyZhEl8s55o+Tg30hqOfWVXbdbWxRHzesZ06Thh9AAJpl0INZJc1
xfiQao4ZqdqyRz8qdGZ6YTxruo+l1WTmxk7kMde4O3gRoQAV2sg8UOndN0vkQdzd9hxvLFyOBz6w
Ovlq9GyBhehWMk0hDHb/wBh5DQMy3FR9+evkECusu4eFsh4iSI24Jw+dRZZ3PiLHTD1Q56bTdrZj
KnUorojxEb+LainHPsPHE+q5FYQIUtDizwv7Wne0Xm2f7pyefXsT/qW2dnlTIaAXivQc8k0nmQz+
AxJgbvMjvWkbwa7g/RY3UMo9M0drqQrMX0QG7PP66GB8mKEuaKumLS2+bJfB0wwyc4SvJPteZ81Q
sRZWl6Kgawis5pR1ByoaBZzsp7yzx6GYbvcOn9kTZt6hi30Go1w/0OHGpTxcCxaifQoUKh5oKGGT
6wqiVqYbzNgmu06bl00SCEVRN6x7o7m7ZpDvnYkecazTr2hxmwn3FqgQH6VFDwgGvk5PWP1B7OGC
G1ly7WUeYBfugboC1RK+Guxd6i8rrVfTnaAL4akD0/tCUwVIphyEHBmDNQ8dc0mDRSmdzpoaRIp2
gr/B8EgDNu0uMGJf+Kt/Ls33jigiDC60ErfiHuGkfmIql1TQ69YaGo57Ihd+CIkBBRNj05mpy1+y
sqHWLUsSXHnLnKX1F5yOaId0nqKjq6KNJmCUC+Ss7ExugGHGT0WvcayyKVgI/o2qlto03LYqidp2
oDE+ZEFzKG09jVi8+zu6uI3cRfKM2lmuLKw9VMdqV7aPi9xav9j/y3ftpT/N+SvWIRdXGEx4uh6I
g/UjeLjilBZvzCJy9yv2IQSWyZaiQ1WIDt2Xq1WUgI38v/eQrPYE8E49bjoL9L3GQzURqaY6Er5G
vzFsh1FpjN6xb8Dy8G48lFQwNd4zp7tmDcY9vuO5YiJV2rceXBh64j/dAcuQ+rWp3U/uOB0+p+lR
ZifJvJAVC+BmJ0vjCEeTGhx6gLagxHwoOQbcUbiTNgLoB34gRKDadXHE8DPVgA7LvtfBu17sHQ4z
Cm9mrRGranGDy9aMZ5tLXFVse/dLTtAb5trrJBU5wGIZnTh9Jdc3H4enZP5SPttRae7rum0CApO1
nDqzQ5tEhrAefmy8E5MYOcEJhSm8S79oJlpzbtiTK4z0EclPsELzVxKCi4tE8sR4G033FOV2BsTh
o/6zRJVGqxEU5hkXSvJfyn+Pk28CIp0NUNab9sHnGu7dbnNHepWiVGhV9y8Po6tvTiYpTiXuh1Ei
QVPyTa/3WUb7l5lXouh+bCubq+CQyxteaKQlbFAqgcX5D3xiBIiX0YnuOnQ/a4Kc2dMgRAN1blDD
CbP0e8nc/hto7s3xP330hJrv31kHHphVHJF7d2f6gYPB7VPCENKKxZOsZA67elHIm6UAJWB4cbzl
fp7jHyta42YlaiWUA3IilTt1HanBlnW2pLZHv6dONMqL0IFlvNRpDFeSru4kgTVskuWbOLrQQHb4
PY3M8T76b2o9+SK9nBxveisk4IhVCRAPF75333aw7JJgYY6ie57DlUh/ImrWTwPehWNx0hRReMFs
i8fxkIJU/zCfJiDg+aQT5NkWsN3jCPriZ4J/j6ky0vxZgY9YDJI/y0uYZCcNOr5RWSLzke487akx
bUqlKp1cXg4sigvvgS6wXOcMN94T4whDCuPtg2aUBF0yy9n5eIwi6kFkEoNHw4EvheFNKOEWEUX/
9yt9ajWsEUAeeqfOpjS5AsNGgMl64ce6VqNsjxmdTWV5/jqO4HvgKV29RR4QYxGfDEgWdM/wELW5
7c/ojTlMbH4QrLghOckGlI1Yo8HOglg4SErOtK9CO7PyyEPSNhk89plELIZNYxC918B9AMLayD/M
7mPLqTQRJPeKS9bK57JLyG2mgHoerc/8TOyajV6166Y8qo00un6rioqatOVrQwka66sePXkIPlcQ
sj1DIZ44IJmMi1ay5EM5ntnlHCEsEYV/5+xiWMpoEeO7Qyq2Tlb8t6iT724wETQlFgtzsstW5OlI
dPSuTl+Nx4Y3055vTJEEOBlhDTBD5aS9Vsw0ZW7OoaVNfTZyqjpBxqYD+s27VfeWZvQV0kYp6lt8
T6q6UNU9DineXqETkt0me01/fgECUuDQb8W0If6bYt6fEyRK9AgePPleNsnAIDHJjOjS4KqBzKcL
VwJUq3PxM8B9GZsvkTvXDxWcaUT316iZzhzywx2Lj/mWRQiRrtZqErO5Rs+wolb5YZ5RtJ3j89rU
IGsx5WjW5XpyhcJhskyZH3wOcsgn9o9dDRyOuZpFmIOrozHQjm/W2fzIyYPYU9vOhcrgxujE3CJF
3/dpVR3kccXYuFq0gcRtm7eyaIkhqX9+rax6LfNEs5Cu/lkEI5V/8z3MfBKfIsbbzD0UKUTomsdm
JFouCmKzH2KsAUDqYIIDXFMiHfABHOeFQLSN5mlaTwYrFNbakTBCnLb5qfcJagEZXJQuE15kF+gK
4GlV5YEGdmdkAew3ZtYwpnn4aJpWGOOAPx+FHJeBdAwNYosXhw7YC+5QJARRPEFJVbaAboTpGOoB
dpwkm92S/bP+19dfm3h63n47FwA/Ex23LridFybRYyFUraLgxRccmDmpNdrH4xDSfKH3N1FZ5JZR
d6jq+0sIBf3VYiGYE4GgT4AM99c2B15I7MbzxtbGaZzjnAG2Iv47EQtwMfaONUmRxHqFBSYm1dZB
iqQCYLU+onAy6qJhE+BgM+bFPkjsKsEvcrxfVK4DyJ6FCnUr0z2nRcDV6ccc5fLwNq6tbx7Cbimg
Rj066tPvbTVpEgJY/o6AItu0mCAsLhtrXE1u5WOYFjrUiK0/ACV+sXK+mrzpCZyOMztPyPArmEfV
Ljjxq0p4+ywDEEgrkP0ECIFd53qBO5tUD3ZzRRkV6oqajyneTh4+gQdYqmmIKYzGvqv6ps+/+yqh
RXZ9DisUOk/4+3Ko6dRD0Gbk4FLTfUe1qGH5SwNqAz4wZ2IKrtrZ/D/ir55yqDDkO0PVAH+ZxGJ7
Sh94edPlrI4Mf8Vj2xgXH0CxtRzQF1uES/rAWYUaczIXNNE7NgBFQMtRsxlxTj2up+a3wtGxn2Al
vGl8ggtTunCIdObLX+U/aiyOiqjfbKRyuRLOwoTm8yWtGeTgqpZspmlST1U/z2N6+5PPHcxzbWP1
FejKnMXrLpK/wPFsrrcrBIBPfURNbq3KaKEHNmnPBfLMY2f2JlKYhTPfitHVfgUH2Rrbwm9SPeAM
XM3xG2PvD+buhw1/uJhQKFWebxcutF4HfAmUzCjBDwOjq/8sBCO1lXiFQ3N794Q62oo3Fa9o1fJB
qKpaVc9DYwFYv5EwxVQcjbDxIf13Aq4mCKi/CXT+yuFc3q4uiQO2cgpTgaxXhchkw+8apIZSaMG3
VjDddYQgLjSt4gGfJnHqM7MMvfavoaqUgPtm5hhFKD7IT2t7tRHSC85KOqmwFEr1DwQKduMFRYDV
+1OCXge0sPEv/7MWfyOZCUWZSqW5lWMzo+pvT29e/cUfED9Mq01x5jFAFXAI1q21J+uG/FteeEYx
k57jkcXGV8tRkvEEAqagRZlFcirrO0oYIm8/m7kPadwYdjBQY8OL2wmPVMWhz41h158c/UyZAKL5
J8AJNFpCHGRtdiw3voP9FsBD9k3kidwaHpdt2elzYQU8EIj5WBNaK9J1iyPtK9pbUaDTkyNKWlhq
k8PvP83FfG7Esh9kGxnmY/qxy1qeOKKcLZMXjFNdbtdeS1XPTpHwkPrwR96CQMp0n3ZbHy8+8R4m
WCr3vqyLdagfeGeMU5m3Ve0o2pnoBUVX6cp2e48IgGK92kIDxOvddzlIV5fYSnJgWwCn1CyITezz
8mV475F3yb97IQqQBuIp7H/Y3eWA2OfSXFCSiPn/GEsxe7mtjos10Oc+vAsbBhZ/f34odb70iimx
MwqzmyOVx7CYWJ74IPRmaaCbbAnM6uOtTVMqMn51Ja4dkydT20RzVozgrw5vTbNx06bfgb6dXKMT
qQi3o6AAiS4cIoFZoP8Fa0to6W++YGQdYC4dHnvYGkN4dMgX9vkVvc7BnopEKmPPwnAtb//6vCtF
KKF978/odnjL+VR00SqnomL57vfVXQwYYaNrRbPqBbVDvutg1Zm1fbIX9SR/+nKVS6C5rrs3dE3w
J8ffDC3KutCAAllkZANeIoGc/1uSTSfRO1pvnSuwCFw4GAqzHaMrCOJmAS+r3x7VJhJjQ8i1PRSh
SZlxQCxZKiDs9LY4jx1RMuQaC1dRkQJ1iYcc9oiUOVW7FHXJBIkPxmUnclgj8ruovmf8pScM2qn+
9Wq9FI9AzA7RXODZZ8n4wTNYFxEWalFfZoSaxhfk9oCoSU07e5jfMKQm6UJ6KQHNs6Wudv69KGvL
JeX537RRi/3b4qwvziEtPjPbGCU9VolI31ZR3g1gbjnwRPMXWDt+i7A7OOBJ/Z6FrQkaKkwgqd7H
NuCtTIlVjH1FZqCHyDpXNo0OHbXRsXZbDNlFvjY1DhoG3uGMEUQhurC/ygejzbbw+985R6FCp27s
o2dzQFMMBgnN9zxFo3yDXCmzl9E4cHJMJIGGcjiQ1sn6w1odfcGReuEyIbKVlXbv1f6Ivxwxm/io
ismh81xHLO8mP/ZC4nXRk+XPODwHSPC45/V8S2bh9eZZcj4yzO79cY4Ixkfl+eodvprXybAMg3We
2Wsnvuganl58ayAMXAgZVL1VA2Y24tl5LmV7Tv8P5Qu3zVcTz6WZWuWcaUoooggQSxF9Z/9B/cZo
MEApUe2qiZ7tcHlh5MD6ZD3YFvnsA4cOtowaj3yAT1WjIn5gf+nBUOj4pLAgBZrMOcJx8JlP3A7r
zzG5JaCSWZz49Xr+yg6uXvvu7yVe7pkQv+eAwIx3oxuUp2Okdu/ghz2LRVjKCjcFACG2RqG44b9j
aJQsWgsr+csnSbwZj4ZMTK1mkqvNoZzljwsGMAMxyZbc6UEgbVCZm/ymK2S/IjWEksHO/VRxd7sL
gWsUdXG+WtE9z/ssXYYdCm+xDmPm4PFHgI6GRZ3Z04Ndq26xlF7aSX+Y5iPj43JqRXgd5KjoU0x+
Nw61ptPCuVLBLhkYqjl6qfpuLXJaAt2+tCMLSQ71jqn6mUlzpanCin53e0pyqgdiCbGYybEw+qXn
29u2TYnMdrn77aONnuKqA1Dz3Y8QKZsc1REO02roBQfYynaWhXF520CGYkfawS+AKpRCxcz31KcL
8DGvLkaKk6Jt9o1/lEUI+GPWqDUjtPb8CK+4g1E9N2phZtmb8DG7UMKnlNlcmXIaKx1TbADnY7rd
HCsGIldbWVA+KbxQDT2tWQR4LX0hh5bIiD2U4NLdgMwDj5I5iw9Tbo1bx5MN55MNfZoGGTIeNM0F
Q7Jxjq2n0yaLldpLTG09607OaXeSyLEUx3NUf5MNq0ZcvoOAwVjHSJpc9j94ddaW97+R9td11rNK
+6KMFwbO3/pO7YSAENoaRX6F7gCA9BVTsWM1H1mgQLDk82mT3626A0gLgbm+uonFSw8shqcF4q4u
RM8RZk9ombvn/9aTh4To5sRupazY3LOr3mcU0YYoCktQxLEK6mxQDlYBbjXZN2AS3zaZGwvZra6E
ENysh/Pjl44eUgIAA9fgvvVs1DAulP23QFmB55fq14XdjYVI9YhiYtMS+6ZTuViWnEv0IwK2HSTt
iFS0XGh2cRMyZEUwUvuhk7Uf6FubZh3AZAy1YLB04q3X3FO29dgwIsDr49X7Xu8Z2qv+VYLra3lr
zb2w+ShD6nHfSmxpGxmaQqr2DIC1wTIDOjgYiArgtwZJzOcyDlZcNgN9JLpX4ckjsgrWDaD6ElXy
MXCKcXlcVbL6LC3araRPoMM+Uv3ExFaJTjXnGezE+ASrvYGLfs3u5pAY1i/H9rLgOe3d8IZJcJXQ
OlE1sWzUjUNugXRoDTknrLoWvccwdZNKevbxAXnXPxjs8YpWP35gveYXSaDPJ4PxkHdB5kI3IcfY
ITymj3c5BBQTZUpZFSzwLTrH38eVBy93qZhk3QpzU9Umf9npRzeCBxzcJA0Td7teRELrsMlpJn6H
aokDKkRQNwtaMsStJxQhDYYYDHnCKEe1ur0j4mEplaXH1zOAdmMYqaNyE8d48TcUXppqA9SGs96Y
h8qVZKmX3NQddtVlphX8+6W2jhBul17IReHXeLN34dEQ9V5CQihe9jSHux+0T31xQwc2eL7ZQESf
5TsdgFuoyZpVAotEPdB8lwcaKxvWRIsHYAiHYgy/GRu0CJwy+TKuZZL6IwgfFMn1YTISyCOLJE86
ubYmI3gLhUFLplhmFWffztKIPa8t/BhFO9UQtihgOw7/h+jxHr22pPCs4Nq6HbSY5caKHgdhGyFO
5furdI3gyLjgEHPgcTDkUfgYhsTnGShfWEBRSq8Shr7MN0LDoysCg2T30ZnbTUhlOpTV7p66BecB
0fyfp7lrGI92KuigBnrYeO2P+vv3jevTafjkAY0+C+8ijDYO9bEkoE3YvG7A5pApu3qSJQQEUgVg
E+4wIUYu/cXLuIGez6EEkwTNtfOKsjS9PFQWB1kRXdpjbC9xKlg1N1phQlI9SQ7rvGradrEk1RGh
1aQSBaV2W0vYyyeNllwDI/arVedMRa/JgoX5Dg7CrlgOa5kRg6iD/yOH5kJfEfMcfzNx+GGyTMK4
AhD/0J3PrLiVdnIj5WA/zfDBJ8FTTznlOGA8oq7Y+af3HPUzKMlWgmkSbOfBTZI3BmSsWd0HprrF
qMywSjIuT/eE1PW8I9QW4HeGwitow3kUI965b95fd+hMMS4vkSUq+7WUx58a3zi1vc/iAVmh+LCH
fmH7O9n6zfg4TDO0Nz+mkpSARZT541raFJwEiiE9Do2UiIdGKRABjbEtzMl7302FgjhKSdiI3raD
+jIlBKgWMsi072ehINIMMbrfG80nW61dMkM1aUE86QQfYvM92jWiihH0Wuy2G08zQ7MyP4U8L2qS
IDupMz2QI4BBTTu6vKm1/Jeh6QdwLsJzGBNuUsJt4b5yddrcBdPSbABEDR/VtQHA7t6QJltaVfHf
5Vj0bdHHxiIeGnkeaAEfJjccaa5UYe0E5ZeEH7DI9IawQZkVf2po+yMQpxVLouobx2+tFP84t7SU
vjY9+J2tUXflv2pp51v5wbqBymA055SWgEg15T0G1dAZQr6kVUXNSlaVjKVxZ7VqzvyXGR2iZ7ej
5DPKtZGWGNF9UlelrTqfLdpRRnu2rIxrv1G9JUgq8JWQ8m7RtkQPtnqLkDB9ixiqMsvoVL3+CNd1
EK0xh2g9R0HKP0HSF0Tmgdzt7sXCUQrz1vOrgpEwCNA/uFNXQKorbRwaOAhGPo31p0rAKWhUhc9m
x90HYsX7j7DbASdCO6mumuy2TF2Mb0EEhdxS0mC16Cmz7UJvh/AT45xnSyQIqAQ1E3TR2g3RfRIX
KdRbaLXlF1wNGeZ5/CwqxaXS4jwJ5U4RB2sDy8yOCJIH96fMqZbecO4YTex8RM4kHnoU7HqYYE2i
0fIiEGNsqhwY8qxyyXeaNmCOaOXGTl2NPrRxC/QXa9+wf0Zid1vcxy4S/Q1n8mB4Ymzx8NslDjNJ
atHx0oJvD6tMycu8G+KSfQpNab7oFGPjwA0+j6itUfdi3sQjljVr9kM6NfdpxlVAQS0WN8RXdtFc
hk2X8Ek3WaEb0CLVQ0DWa0FxiXGB7icsOWxJ9NrZbSSiqpmgD/GPavaPdujnIYyU0MpxRbnTgh7w
Ga3jLMCgCLmtx1c4oMawyN8buGpTQoU+sx0WdgS1jUimeTnllB6Mwt3YJPjvskbqWAWbkPxFoYgD
km2pKUThbG2LMtAZJUd8XeSdkVWjV4tJCjEbMA9E4fh68hbnw+kMNCYPblb+gOWOcaAHQJW7OI2J
X/YxGk6PJgcjqj6GH88wDAU0tKRB3zh9i2RE8+gzp43vHRgyqW5yw7hKdls8TBfDjgIeouZSgo2w
qV6PxcVerEOYFLhZtG12eBUBfNInUHyHbh94o1YfTwPkthlvnpHu7cmtuaZ2kqja9Y+J9FUX9Lh/
o//I1K0dcwwpvg2iX/Ozyzka5tzhzTo8kVlLO8EjV11BdHBWw0E4gdHv+fL2fPzRfTZ+NX4U0SX5
MRfe6U6M43suYKBpGW+EU6H0hAPU0v6s+NqyRtOWREooY6MJciQZDBz/4xHESq4MORSrAU6LEVxL
UAM4wwJiI0PCpqkJDdZa5/Fx+1U3LGOP0aDtP+6+3+0QD2+snFJZ/fTsLh5MlZMQFMYr53wg1ade
N9vgD4vjEBAoN3gO4XMymM7/LnuD2INSq3ISAiq0NJtT4G/Lbgf1ntEJRXXBlBkvQEOsgkx8bADe
uYdgUAWs/OxWZ1/7t98MTCGCxnsqNNBfBvJALTFGT0ZILO/EEGYUv8M8x2GwgzVFTX19i5jMBdlM
fLqu8pYXcUOcL4b/AvJusZ7f/09L6fYrdx+73QpBO0+WvaHCD4BDtXWwPxJ7QdIrdmNXg077/+1B
Omco4PEdcaOtmjkcotLvEi/A0wE1U9SNw96qMy7VCzyfWf5hScDhAQnQFIRbBcR9CNGWUKh714i2
QVnVcVhHUfQoolvSUML6a8cX0WghDNEmontzcBoaWiFerW0NcBzmCCZoTIh58kSYTpduGMv93M0B
djZH3N3Yxj0+R9jopCOJETTEff8Ls0vIwvS7MBIsBORodbhpgtiVJ1/wMkQR47lFEMBql4X2he7j
+vgQlgdp2tIhCjBU0BrmY6TZUhuiTi/mT0fgF/Mz09BJkVq5SeHOLCR/nFUZE3hKDg3tmdgdT1q5
qy9lm2u8Ex3VNDJMMpot6dKDtpkmZM33Ul+Z2fWgmjSYwr5Cle7XItnTiqOvEavpTv7rncbFtlUo
0NHIDrEu36s3+BIAoQZCJvqtuu8NYofjl1GcSu5irCxjsqxDGC85N1RKSRmyo7D/Pp8rJeVLekY4
IH23jIEjxa39w4BBEH9mBKf7rT/pY59x2SkZJGOVx/x/4aZVc0NdW2/yG9MShqk1KsEEKfP3+iAM
AVU+t5qi6dDUobq/CJRkFPsrrHgAGP9yRGHD27NPgaxPL2yyG4gzW+5bZ5jnup89fZFVEqYOwLGk
uvtU2BQIte/jNrXpsCkofZAVdz3YyTD9+G50Z3m4vtqadRbRicGjHZ44A1DiimYN5v6mzvEW8zip
b35CnM5ZZi0Mr/xIMUUbBiWe2OJf+VOFd3H3fTQ/6CsURIN7QB+9fhO1U9y4qn7jpD6AJNcOL+IM
cn7nq9Bmj3au6yRme3G6lJwOPXx84ClrqSjjWDpNudM8aWW7x+DwUEDmWl44DJ17WsX8+BDawurC
FG+ay03Ok5HNtmnGwphkUXX/AyZWZKvs9LQxh6RQbk+uy5VW31Ct35P+BM1benWNBuOSOAXnTeyQ
XATZl2fxb37xw71CE1HTRAhILlD4t8mIROhAo6cfsAy+PfMndj8nryEpNJv8QTfFn+hMy7AEDAd9
fIdt8Qz+n1WncuSWtzdo7b7DTTZ4lTkOszOt5Ti7dRaGOwfD2b900UUdNupft9bEviCyYsJhZV6G
VYsOwHjw5+YGREKrmItHF5HjobNxo4vVbQ1R0L3lbqKTDCmfGY23ziy3ICx4Wam3Q2tdQcSJOjTG
BnOQGBvWkMlvrvai+2HcYnlUsmoY9UwwKxR3PlscW99B4/RlbkzEwUoJwM60t7Ri7nAqt+7pGKjL
TPQQ1PoRdvJpq6L7IaE0JT4zzK8/GbfzFJsVJDCHjWMwLrXf1NkUcM5T66wRXuqMFf96HxtVkqNN
Gwz+zz3t6HbsfOIc812LuM2t/pp4hxoJWSdL90HyQiJf5Dxb9AiNLRh/1NYa2X1JD40LEHjS3rCp
fsPFskg5aqdArWom63xPxPXTpP03fl7zr+e8NdJMQWLtDkllEM4P0VENJQPo7cGMWu/zGbG4zBUt
8DoJ+lapVh1eh8ilu2SRUsDj1ibsewQW2IcxGmaG0B/yAT55meUmKcuNSNchbsdzTWV4ewIpP2iE
iWGFn3pxrr2xYpNKR5cbxKFKq5Gedn0zRw2vhWG64+ZrQnyVCinz/pwe2GYj43xFlDWUvEisrEFI
XNpfFYKqtePQlIShxIRgW35R+sWpXySE5F6/COgkZaDd7wqjMRBdo4P6wv6acpgAV6wBfLvvVf3O
qHS6X5xNETxO9EDpf3V1ikw0RunJ2R5ZHuSkRDzc3YYM7MnP5KKwHSgOpE91rvhC2kDwDZAn990C
yoDVP2XVFawLFo3NEDyvZoEdHqDUiQojrac1oo/I1lSVMEr2bhg2wVPZC+Bqomw7pDCVcjUdIdRT
cQyI4Bee0KzTvcLwk0RRxklxp9fAixXgDPesCNWlqLOFYu2dS5VxEuO0pLmnsfqf0CrZuBin77CI
T4UUguMcEMrHNNTw0FLXXt7mL1sIRVYoSlKhT39wbpWzNUg7QwjQOU/3jmBTyrjyw20Mg04Cs8UH
1oMlXaUbrEVpfIVYw6fzDxVTm8vZwgQxJNDPLTOHr4OVnaeV5PVJqWD9eTO2PQERpnDMJ81ThQDd
Y+k1XloeBbwEEUtSQSBHhW9pWVogs5wqaeFyLMTKn2BinyGxlTDWamzF49KQqTBewVr9Uyho1ldI
6YV3S0NcGPH25f234hysadLNJIUwMjvd3KJ6baB9clN0O4vBKocRw98OyBF5pq5U4o53mZjl5h5s
NXvqY48lnfz2F5a/3C0mUh2+s2HjHvSN62GJhAqfHHGO6OlqOhrqkJom2hVyugwj7+dRdd2/z4q8
wY2Q1l3SSNJFnxUhrcdoCEaty/ABA1R/wy6yI0cGiE5BueZzgjzIG/p9RWWGPM6KWFCb0Osdppti
nSjrl2XfsBexf2AT7t6slmYMxVoS7rfNCRaeCrcP6Y7Gb97Edy4BRLplZrpDh2yigilND8UpgBlW
91JdoYc/bJ8ZSbx0McVwRQdJ0w0/Xjsdt/rB0zMtS0SdCnsdM52M45qjuPpwsQJdDYpiNZT4R8bb
gBDSYQ0zU4vm02yRlsJm45HzY9nfSRs53NN0ZTa0VHmLcaWWqABJSAe3kox8WPigJAhfX/6aV0YP
9x6p4OgzoD6gafLGWB6tqX6HYa2RqFODIan7Z1VX5NhOumbcXx695KyFhqwY7xPEEg9fXmTON+gG
//qS6GPvPIB9rkjlFOn3jqrcjpvkPwTUYS9Uno5bB4/SZ9o6p87obfV8sW6GmLrvdU90+TqTvQ4d
KuCtj9g3rjnMv95WvAs3fKAniImijQAZK80azJIpLQtrJhbzSRa9cJW1g0ggKJywcIEVEfVG+UU5
0zNftcsl4T0TLrXBpvyZ0gEbwjbe5RTNHldzFwi4eDBeLTD5fzz6WpJssyQUY2vOcx0Bv/43fdrz
LpXNjM3Muua8j8TKkmAVBXIOiEPZIlhpJKQwI4OiNt2mNu6n2/1yJYnP6h2jDgU6C/UQmtax09Ty
4MI5t5RfFtL9ZZusvTWhWTp9wIfG23Zs5JdzRvH/gNd0p4neDejsCFHbteDbI9aWtX5/phvXi3oI
iYl9aWECCvrOHn+ZMggXnZupE78n+QX4Ma3UyYpDfmPJEPD5LsYv7RqZI11lVPbFW+7VZDShhw9x
GNxcIIAdlbOGnhT39Ei8nI7GVgGl5aj3X6SQlToxXKsm88RnZt0MWTxW2K7ttvxn02wnIz2+Gy0R
RpbNWiw2h77U/l3J0WhAnuIuACR45dLHaa/2dhztDjdJCCis/mXPRD8SOgl46GKuAsc1WhFe8U+e
A5tRokwTm7edHLjk0dwMhF7l4MM5ogsMG8Yvgx1JOjIJ4peMqIhLopelyMxSkMumy4FYt+lcIikJ
OU42qsJSs15/iiESf58rap3Yt0vvJH893jSJL2JJgH7jsTawP/w5frlo8mMDnlYlgXfwjRkQvDnC
V84fZsXt70yT+UDkKd4enGlcXJIzbwD569jKwPW/YAfG1irIYIDkdq0BXPrYs2TviSTWedUpqkbU
ZIke3SApquOw6D1okjdintWhYHz24tsj6WxNbpVv53l3iX21enZ9+Fp2K12HQrkoXXH8yrnMWFJw
O4O315XL3iRYJruWwwZ/Oj+ntV1QCOSczYxb/8kGIDdFIo0xox0hG4bvA8ZzlzpcHFDuYOGDMSsd
D7PtTFG4FqHa9y8JdqH2OHQqAFChMptl8vyocv3CuMtS/5VDhegQXryXYfg7e4o6rJ2rI2cfr5qt
bqy093WUf5xqDGGczylqbqBAraX5TyvPUyviO/4FrkM3Q7TtJwJA+XeB9ngnr+fbyN2WtWGtj87Y
qrmFoXY//FEuDwUhi7Vh2M5A/fMN9EbCsX5Im+VKSkjDSIJtDi0QwEdyoAB5CxxIQggXW2UF0UM5
hrLmyx+jIFFeHV257yI8YD6Ft7aNlAKX1nuvXZzAmPHH/SOib4NAA/DsGwmjrStdOv0J+Ha62qq9
qb893yLvPKUPH8nQt6epYsmMgXcYm2847AxfyjxqJuKPbiQMDvHiSwelYuAwsv+YGZSg+JbTSsIh
4b3HQw+JbOsWKok2vRcTsvRMiBsnknX8GpwV6aD0g5fcJbLPMdqIv7e+xAIBLypVanrDpRkqKJOw
WN4UGjgCelNwVjO+WUZ2aX18f5+WFYHZmWMAIkfbs0xkQ9Dtil+KOY/UnorGQBukKoplaceK+4GQ
hy9UtyWW78Mxa41pe4/BXLqfAzv5twFmNKTI5tMNEfmmOjgbVLBKw771cF2ztYNVfSSLxKF//bkV
VnpFbkmnjY4eHO5LlP2cUSicLoNLTopI8ko8JyyOigU/6yn/JyWj2peGwt6m/FO+wTRgr+3OFQ/h
UXDMYCgB89F4cANxDovxcGxCxl0HEgzK/5a3f1Ic0kK7oXdv6U7LgOWuq39UK708N7PuBAEZgdaA
C85HGqD6zoUhPhlIZ7r2Nttt/n9G8KhjSgdre+kITZjClbUnvUXclCMDrBxpd39TUxrbKOad8Raw
BMyOdkUlD+cisrz+DVpghfsKp0kLUihERk5+Pp1/zKPU4Sj1ccu158OEYRLTHviig8gLR8+m69Np
Bw7jDIfBFYNU8GZxA6uOTHN+cUSTOpWSZ2HAzBEK7E2DY83EXXO/xpir1RNDSM/dsvkXf72/uHRa
bVidaxY2Mk9r/HVzSvlzcupkfCt/aSE0d8Z5dESQ0PG+wzPK/zNqwz8K0pF3ifKC5g38QFSwr4mx
NN2pvjP85l2lZB+0MojjhoKXKnlokMuHM8P+f6KJRrLVebilD0pI8VDob/DvY1RsjVNUcqcDKY9+
6jJFC5f08569CXkjyIfOuzE11NQd5ZJDLizi9VQJ4OFYHBOltLGxZtUoBTFRyrl3KlzL1IuQLu9G
HBcHrowg1YrBCcyD40/wLCNFugOjbsIUbkcqCKhClu+vcq7PGPc5mbyj0E0HvdYcfrDwN+mEd2mR
ND+JCv17t0VjUZIvJpBPNNqy/fmfLAuwgvUSkF0NJw74n3Gx5v4d+IRMDujXz6tIMOVLWe1ad35h
D273couFHbX8rD5w68qzRc1tN+sAZWTnnjegBS14NO44Lxqw32w0AtwJtXMe9Qr8Pz3sg0DquAjy
hBunCl5UPq5Zn9i6hf4TNvlA21ozAYFs1kF5L1T3ZgvlIyL6ApYNvTbce2tZcEWoIqbnMvgGdSpy
yP2ZKZPOE0BH0KmwxmI7xaik37jwr3RgLJoqBqtrZUIIqvoIWi68/DFvhwpEMMCbvdcYQL0bE7vR
PDqc7/hrwWJDRkSD9dtQ8aci55VvpcmluNiAckfM1SezPRidFkbOYFCLiHCQczKIVWyN+BO7XQUN
EHzq+aR9S6qATN51FtUd4bv8s83NsPcNL95mWLB9wnMNkvUJwDbOGMv3K0fF5NHTQ1YbTTZpWAfk
zDnLI7OuNPPNprH1VYCbrb6IgZO9bqno7z2WgYKgUa8i6yrXfHXfyjfdY4rH1Jc2hnCYWSAkzj8D
tJsz2xG3OJzHtF/45kP2fRIg22xZEcyT094SaTlGQw4HXqj3F8kvs/zb9322vomKBguhm+WeevJP
YSq9XlMZwtkL+WdTovs0XF0tXDXhadtrfyq9dCCNCRwzvOx1HSklPbFCPPIXlQi6YxphRCSd2nv/
bX30T5Y4rg3AaROKahkiPAdcauIi60i3xdEriDKaWOVqmY1bxiyo75un6rcyjlG7WDMJWhQnX+GR
PgsLu0k/i8paj2Hu01XeJWdOa4U19Dpz/vE/DQ0ASABnwZplY7ZGlxyjt3OIxN3HlIE/oGT15dkI
nrOEcoIyGR85fYLWA60qMqedhq8lc84kctokTynRaRZe4juJl+J0L/ZUNrl6GZx5OmpsTnCmboq9
5ZWQA/C0uKmxtW+vxetg28wBkEs503zCWZSAwob/cnduYZ9e0/l2v48UQL7ACy7L+2lsdGpNac7m
1DJa1+FBRN4Rf9RBnBgcNWZFdsvNa6WVwFLGf/SEflWAXWJD3WfTdzaeZX1Ay16QMuOy18WDRTV0
R7y9VHwdS/sE4GCNWIaX9yQYIwMfMldxKQleTnOSUZUSHmMv78t4KRtlXFwn2+VL+UD+yBk6x0yc
hwphBQQCkPjw3oqXfr3s4X8a4rfdMeYNswQNesKw+aHHfgu/NqsgZKbtF4Q33r36yeHGPciHsiEf
KrJdnx/9rMWSRxsNRUKqEEEsIbxYVURtzqTQ9/VDMJ7sjwUIJtTcglV07qaLIti5lU2p5iNuWWAk
MudrBvIA98PMq7SVOrfStASlhHfdfxt+sFnegFnogqAqbx0wtOBEDiazPLQsKjsUcyDpWO1XcHhv
+3N0RUrWHBaEOoLTjl+0txk81mz0rjXLkqVsyJ34yRgjOnF0U/2jrO+/6M506AyYTc7Mb24c9mxw
Vk9hgRHGx3/ENBpiv/4qR1LpUw8mgg9UTCgVGnk4jurucT/zJHcHn/wWTozal81A0lAqfiJe0AH8
62oy9r25d1tiHrNd/MfsfnpzAUfNlnAlIhP36phgHMQB6LlfKuqe2AiaXARF5srSo4dek0OD/wwz
fG/C8TiNIdFxpebnTb7aOXCVy/URGJEtXzEtdUi2rjRA/o/e5CJ2RYb9qF71puemVL+QVHNzddci
eEVhEpOxo13uR0HZHtKUo8cg7qjuFNuntPXJfvXN6cor82nLpHWyzpQEZ17j1zJEQkaQNewSCnOW
gWuWOM2k7bagHaGEmIw1uxfdKXQdmSDEz7NDofHP7lIGrLuBiDcKcUDjiFuUlB91Tt1QOL6mSs1N
Dz6XZXnJp0nFtrg+60fP/kLLB8FmpGF1l1TJuvlPEM9PgUIsEX2kJkJxwjc7w44qYi3qpoX8xIuE
YvHbgZNOS4fQixMgY8j4CGjsDYrtJL0b2msoK5eXLwwmH969CnZ8KPA8rA2SD55G6poijxK3Eaq3
8J6lS+GvjBQB9dgyj5p+BtuzPXbLY4ecjizQ2igcGNGrFHPfAjy2OP85pzM2zQFFwk6ETzCuJcon
Q51f2dkZ5+YJe2UB1GxEOEsKPYd2iUE6g1LR4CysZOzrmvYd1KfGplVVsYG/3pj425tVI1kf8tps
8Ym8nARq11d0K3iUBavOsA6TQfJ/1MzT/r6Y2XSOXp5Hy34XhNWI8hGIcITSzMwgtUGwrZkDYcOL
aroihWsk79GTSBfhdnr/wV8Jtimt/SJXycQmsB4tYNa1D9P1AU/9igbwv55yEMESfW54eVBCJC4h
9zm2VQpxDeBwJP8Aal16f7OjtNVu4vkdoVXRKrrKPCpAA3Bv34Z9iFKgn7VsVzR3ayHQKUDVItTl
+EWTfg4F4Z/+5fTX8KE/OlwzkLUU1Xmlca9HSfI32x+9mBzAwaLpAxQ575DaIn6tFKUhLLBoYEzA
TBo5NRYcyRMmRkvssFYus3jtFkaoWj/OYLiFJrwDLD9h1ilCBSuRrCDzYaQHsCcKvCKYpQmy1Xzt
0KmbLaia3fnUsrX+yrwVCbpV+yr1huzwXPXSLZlBq0xizA1gdNGPKqxXpb1rwj2gtLKveopyc6i4
RC+rYsBq39xyePryL6PBW7sp1L8V6zLO9TmM5andRFWYNkdiYIK5ujyGQBA77yMT8OwRUmKfv6G5
7jfXEkg0KxTFjwE6LblPkc9XozgMP5lDCkwjxfQOs8KT0Oa2Y+n7P6g8zDKHH2djhhPcDNdmXoJH
+in6CIWjsJER+I1V1iDkfI159I6owFdFwI9mXPFhLjA3yIvAipDLIAEBxZMuchsgOhUdH4Gs0EiD
1Tn1fx3s4xqEMsskMW0O9ks2nemodiKjUJAqFnDLD0l9KP51jS2jn7iZ5X4pb05JetK4P9dUSQv1
pefbXTjmN9DzZ2oFZJpqPq9GMorI3ac7vz4I8CIqIltE2hDfOw7gdFBFLxkwI383L3nOofhMZ6xE
ejln6iXKDa77nWjzAUm3PwKBaObHRReekhn1kRlyqONxU9spCid6kjQBw2IJ6ENOza0mT7j78g88
zJORMBVi4Ta8oBCxSaSN6ohUwZZNwg3RnY1C2J4+GHnLXOA6VPsHW0AVjiuO3YzzPfJ71mZkE8U/
pUx23JZwE9dNVXDB88U24fDtCXTlvreIMhQqEdKsB+/qmbNdtYZTi9lTPx4OSzH7QtU4VB2Mmm5Z
qPi+zsahy2jWQuCyKfOVOgcSvt5ybGv2lglkXuUAWkP9H80FNct+1lxbYyYoFgM6aa0LeW8//Rsk
CKWmdh7Gu3QO0yyna/wtWTAlVayGiAudUcMMV6WeyMsouWOfoozXtUpPgnaS7L9tL2qf5EmKL0yL
aPayCukfJxEBFc8VnbLUnbNl5ze+pyTtHwfXuQH2eJwHpkl7w4l+vZ9C7Reiv7kmuD1AdJFwsjk4
cDF6vRe58B59LBmRdaWekpoDSY9syB2dlj8+hDJU4WhkCDf6KVZ84zHQjTvQTGBSNCekYPxOLLvk
asFxGxC+2UU+goc2nF/wZ8wh1asQ8F7LwxOGWywhIXqjTdsZKb3Udr0fZs86e28n3VhI9+iZO24E
/3daYSi4tBzZK+9YhS2FNAdylu6HqVYLgSKpORvU+RNdjKSfV67zfddobhnM86pPFeNfXRC87uOn
O1Z+Z965SBF6Jx0myGayS9nC/djfktPgRXdF2PQa1XZROT33/q582U9IaEGdnDqx+cN5ikbnL+VS
2Ys8WuNbQHUOLTEZddeb2jx7B9slDzB6b25ZaOxNWRRSkdplNDGopy1PWsw24HiCEaw7/sFv49vk
HR8Rv62xDI10w6lgweQYsAl4vkfO9maGXnIvfK34mLPy4KwJqaQ88Lh6dMpp0P4yOQRgzwvAToc8
PzgUg8lkuM7o+WR1dm25f1S+liAiBDvNA3CoXrLVkFN65Y1RHKcOZAcwN2Qyf/AcXPmtuwoxj3c8
9RZBElpZP8BDLJfJP6z8ACnszRiWv1OQl8Z3CZzWW32PNeTrpbYse8/XumBdoEI9VwqaLP8wV2k2
MKBozqvBHAi4y/PJCz0grd2Cqm/wesp7ymFnEtYB/RraYY/nh/vHRl1DLvyZYW/7JBS5pW5xj8SB
tnzs/+ePDoCLh7C2ewERFNLzz2hVdXSjnEjyiwp0xUboSyrpURgYo0ZekUJ58yKYWs20OTn2Wq9H
X2otHSvVyXq4KcDf0peHX35D8FJBrHepVA4aaoEiewO0duNivnODKA0/MiXzJ/b5tj0T49/Ej3au
rTjyMRxpZ7Me1qoUD270dfEA8qNHoUVZVAQgqVq4ANta0khgN+idaSMAcJDPKlVRD6oy750r9IkC
BlBQALOET2a/DuoOqwUcKvAIJ0sR7hH41OBuU9/h7rTQ4UnAMPCcfnE3qlKg0PsCxaMfjQnXcWQV
iSz2BwO8wtlSNq8OUJb2Fm0ydMdekEgjoIEhRc1567mUAWMtK+qhPqzA0AYLhTgCshYUivMd55r8
lWWy5t91BMbTN8+LQsCZpOtCenKiQimNtq5C2LZuLNxw4jhFBC/4thmlcDBtopss0m8N8XGsrSXS
42l6BIti8RTvcX8+nmDRbpZRZm0Bgw4CgG0FJvLIl09IdIhQuATTxA+IvFUhkc2r1nh0tLHngfXv
8M/dcJjsFyX2Gc7B6m5y/5voqbh5K+kPFJkZtlQQEZjF4zO+3tL8nDG6vGttf+qU3/rp2aY3LWZU
62Pv411LQcD0J4psf59h0oAG80T6QBNBPW5grcsI33Dnlp7mMU8cy/MRsKGPxjjblKHjEk8KZuof
aeW9FIaCZxkFTjrxWRwGu6XGCgmXtFZrH19AbS7GoA3Jeqjo/vMWbBAWJHpd6NoHFKDn2YtG46AT
7s+T24Fu1IAaMyFC32PvexzQ0t1xbNKtj0RVrGwCXMO8hmi85zXN+LGLirYExMf/5igWz61STDja
18bzFihuUDTcbLO6lv1T5X7GdMEr9BlRBoTeqKIRllLPq15dD+umCRmzi2y7dBjxXr3vIBk6FrkA
tTWv59SHuGCkrFd27SIUcR+o32/bBzhr93iNhOvd/lv2oPA1edk9xAejUwAQ+d9RspojuDcWPM2p
pzhXp3cFA6oj5suAtWu7hV7KObsEul7+oI9oifLRZDuTisI8nFbaHzceVLL/eq1JYdeSZh3Dx0by
ZO4yPj4PgIOJ4xV9dE706ygIwyoVqXNMk0eJ7Tu1CS95yZ7cys+PaUl6YnF69K2yLLCjSuviF4Vn
DkqeJSInexifWcKBjmT1ZfILqyL13nYDB/bPAALow+XXMw2pAd/I6n8926CQm7VmAXXwoWDJQZjF
bWQw3XLU7RvUKGtCynvAcaSc5HlLhWQ1kDnRHrsIFYaGVTkNbNLAoOqAtRajydpzd9uMs3doYa3X
RNoAtcjla68jWMldjSc/U12wRto0QJ17qqNcDc0a/evRH4IC2Y4kFa9Jb3IOyj9iwozZMHbeVgxR
EOASRsQejQzb89gMQP7AI+bimE79ApppUW+p80PMKFn9Yv7qh6paAbGVzWCz6xSCnB1SHibgQGzx
zcfkTL59B8A2Ne6sjVKU/BNTlH6z1ynTp7H9urSAEoAzqAMxWwrrDWD8YxfJLJvO2QPXBTH+Y7dh
R15V6rtZAj3zfU0aPjCYBb99nEiWi07MB+uIlWfGWH5jnOMryLyVx9VEI0zb017pTNGDqqHZybGj
KlGqONMNFjEA8+sLO3mBqNSBuN3LPbxrho04EjbAkkzEEOZW90ikSpNMlsx19wXqvZQpxOozOyg3
gZrRvq/KlsCuzd9aXKUw2sXRltbEHZIgdcYhPco/3tVHi45qUSr1dfmsr2pSTAz199d1y2PMqVgS
eiN/wAQ8aGWhum39iaDWOd7sj4/OEPmnumhoxK7fqLZObhD4XrG6oac30xthBWvUrAtBhCPQmvSO
cAYhvZgPt4kf1vy61GIarmbpSvDtaIuzVWZPwoUQ06MeXpxFy1v0iS1ImbmPZzNOTTF0sJZdiNSd
LqY10jqwJgyb3/0Vkl3bkph4rpt3b95Co0sKKg630LAw52vR5hEQQDZrF64a8X7/7cQlhJUjEEFT
eqvDeDI0aewX6LsxuYQ1bPX4UU9hCdPGXK0tceG73eBWuMxNKyWn2Mpb//QdQoWOy1RWlEn7wO5X
yl0W2pO9TRWCFK4QnDnAJ2R66AHphEkt7gwTwazeOvbN4l+fRaoZUYXwTzb3YGzUalXDDJWHcRvk
avM0SWxAPaEg1DPNhRGxS06G4SBoLgR7BIXkqkqhERpoZkYrTtPhuvSRGcHeb7d9Ad/E1tIs2NDQ
XRsCUjLU4POCabp1DeIbULp/t7dV738rh0vkv3tTd2Tex5Dfqm8th6QhU3enz/rAjrkkcgwQZaIm
dipHVwiiDKCeu7yOfVTy0iQrwEc8lZufYL+Y4QCxwEDTZ3jx323LhDvZMRRlpBT+/OJwQnvrnMQU
Vf99T3xqNH+pLmEFvAVCjdCs1IHcvpNvJsl4ifacLOOH3BZs18Sqgg3nUCWkr6LWnS/GItEzB4P/
2zo1tMse+kinBgNbVZc27nMGWWnqAdxoVFRQMAj1WaNHByqpMNGboVMEwZQ+hE3zXMbS7e/F9Tmd
UDNZMyvTiuJEH+A7/AHPSjxxdLo18RXfc6/qxt32oyBXjNKHvgEKekfqVpWyiIx0jg3uOGZy42Rd
Ltd76o35v05So/M78s3t6xiukM3OR7frp8Z1TnR+VGzU2zWnVxyI0DrklKQFof/xNRBHZTcGFdMi
TeH/UlQHvN0m0z0K64QxnwIHK8KLHmom+02G5H5TLbRl8dy/wxJauexQCTHqcdThz3JZ6kAXwu6C
CWAppRn2qlsngHchd+PpCYVsikgYjnV+FIh1olCz+gdMaiwWJuEPtEPjFp0OPZdoz1diswrdILd1
2ASGgEnX8tqSuSZ4MtCSgVSBKuWUS3FmHfSmKEZBsPCbqAexxjLWXnAhI+gpHmvoRP/rlyuYgUcB
imWwt52hYkOlEIBnjv0gqNO8FFPPdovjJ0+RkcNWfqAEOcQTftGHw7+uCINjc8L7DeR4F7dpp4/4
+/FTtMqdpeJSpitQqG1Rvpfo+nDrlWPsSMH/bXXyocA/nFplgR03KQs8gd32LSvhSRgTw8TNpAS/
FYxX39e9/dkm8Xd3CbiO+CtLxERzNx2SmQFPpuxGKYoI5U0IzI+AvEy5bvuRB0iqi3YVFj8Q6ExH
ZsEM7yvblobrunsIUAQ6puK84y8fIXhLpTySjlgP1hkB4i/4WeBu1WmAui/UXee5y13vV9ecD6+m
yZ9tY1ZV97Ic+qQRdwWQFY/R75ccIi3aSKNw3QZWXmPCXQ3gfeY2Fx22h30cLxWuhfetM5ccYSb8
IIXyDPdlmlgch9/o34jQWof917PBg+SyZK3OpolvuasDmZdfwpQKBnwFyPe/ufnCqmfYfUrV5mZS
EG2uK/8hadCcsBQdeelhJA8zovpMVbfzhd4mnB6QBkizana/D75Y1ZRuAv9Tb/9IKmg7LkPtn+Zv
+0OIO7xo6xpV65KqaBzDF4JHnltnqhugeUb9z0X3xtZXwlfUEQgRfFPtA2E/lIyAJnroFMgt45rV
tY2tJvmKouVMx4DGC2cvXSf5m5D4gER/ouT/wTubKa3IzsQvcZ77TTR19vF4ldbEG72op7TcgYWx
JkrM+5lyh2FZXEKl452ogcKFvp/yO6WxOUKE1SCAJCf2NbbaZ+oWZBQQJy8H0jU3Rg4IlI3WGh86
82EKRMQ+/grTlBedFlOLhMoqcgjy47dsmfw4zzQE68CbI4zMoj0INrmy+mnyDLx2C8PTsC1X2j5E
6SE6vqgKoj0K50yqValyxrQgTgJ1Gi1VBvyWxf4xPE/IgGtsUuMxfF3PsIGwQv0D+2AeDrrW95TF
xyEyI+G5zMXHGIfLeQwRVPhmAw5vj/m4ZW79mwPDgBOTY+8+Vm37aPDtJQa46yqadytMZ4vqsp0o
LFKZdIq0hCvxx5w3TTLFK0/lzm+LktgDLLNTBWDhV32bhK5uATRfvOIAnShy3Q71bXUUMz33WGre
a2gNJYHiKeSjo9CfvwaIJ/5i2fDDe067mBQLERLGvZHWQ8kbbk8kaGFekKGJ2BZZF/XB0R+AuBnv
1PrrjXos80PFYlvLtK2Df8pZt68L+n4bTv9Lfw1H3PyrSJK2YPpsBgxyN62cE8q83OiZAsgA/Py9
InZ5jiGwzmrcF1Hm/BgRFHq380bQJJBAnTi8AQuhow+S1AzLgqsk4cn6eb2SiRVXIDNjkLB9Ap7l
mYpJmK4Hko/lFr4475+kY/yNH99h+mj3uUY+7ZWEPJAbzSWBTdD61s2K8I0Ez+ItOFPhE0yGlM15
t7+RPqIQhRhqk5UsV4CP6CsQlJCaAO4GVSiI9TZDtCgKhZC6Vxkl7bQ9DlkGGisZuF5DhEh5BKGG
89MD6k9KHKzSS40sTMPTXGvoNWPuwLDPCuWW7t3Pl+8uEVtFgDD4O2dmaGFHqkObYqUNyoI1gF9m
q5LQBLs7s7z2y3njmvrIAHk3qKfxt2PiNUvgCEMOeZ21rOmlSMghBj+Xfm2IaiOWcW2DjLgQHo6i
HYkYaWvEbBzlEJYtVy8t2VeQ38FHlUSx3UvnANB8UUvoJ5p1GxEFN/yVMgFil6jnFq+227OHP13Z
2n0Wz6J9MjRZSK0nWXU9E8wMRT6jBHerKlzJDsWhh+C5vK589SpU5SPsWzVL9zmK6R4NgnSGp7Hv
AkA/Ib9p2p8433fsnsE41tnzI5TO8GucAo4s0EcDX8CwOG4oebiU7WDpcsOIoi1M/SoXh8Qp2NvL
42IzEb+ny06pAlPKBBecxy78HAcmX53kZltoLj7c9LlVFuWoWsIXJpp3ttWg5ZowxonLHpnoN1Qg
Rak5C3f3tsdfJJ1EBnXS4rTcUVbm6gimQqkttfkXOiLPxqh/ErP2YitemtGIIfIIlngnFW10cjAY
H9EXIK8ENGE9QILEUxVIBSxBdUfTXlor+HO19Q9cZFq8inz3q59eNIXqwV7HHF7/Ds8F7a1zt3UV
SG/EZtVuWjg+5FE2v7fefF1k/rf1k6HZZa5YiHAbdsG+NGNR0E0w6LkAZPUIQe4fO9mM4Il6HFcX
KI3KoR6K2q6IEaQbrr0q/ce8hoTwDk1fIMZT2h8A38UITlcCQM6HGLZhr9LfmiwS8qvjwj1XUGcy
BA/qZS3DFyN33Avejuh3ZQkhaFKiWl3nOUPAiu99uxOQ9H1TMwurqhna+KdGNfc3KOoYLR1ekCLd
XfS4W+yk9F/YmiCq2g+6hh1jS9UZZwLoSWGmR3QGDy5zZaUgDpwZetbw16t3/hFxCi02fvHTJgu8
gZhrJwcmkYRlAxZsRFTz+ToCnQtsdpUh/hlVbXOOMhsatDNpoMGX9sqm9PakC2O19ZFcP3ap8Vj8
4h7koW8WokEcTFePkYqvlj4fooojXCrq1KLqt78ny0g6kwaZ0tIMbRzviM4mTXbeq1nzEy7GOooQ
mqyYFnLD6XB7lzIGjF9aWhrC/vX6yAsZsyOpakBgT6XalJ1JyyrD4+4sQGX2X8o3Teutq2Em3sxr
TCzlUdxduO9aIG3uVdMNUzDqgzmgaob+aBWvQvGdH4EiQvL8Oy56OB2SdNaQdXv4yWuMUqp1eCkG
HNCNwWJHR/+gr1PbEJZLgcaJgGlpXmupk06+VoRNS9BmTHxmhmff/dNUGuUDQOk9B5qZEB/FQhSk
i2DuO7j5wSCSjV63TCOmnxf72FxJJLWYcVtXGx8kvL1vPrNopxJz0VlGo0xgxv3j6cqTRQ7lhhfS
+opQjRitJ1TyF8w1s2DjWSlt65V87Nh5fZhwYECHuLMGjdTXVGZKtBLfOkmmiVzk8wCmOGC1i5RX
ob3yGxpQ5lYIeKFyQxXhHt25CWe+a1eyhTVl36GYDG8DqE1ivH8jzvBAsZ+Lp7zDgpTPW5D7CPb1
m11R6YmJ6aY43LOG9I89ogkbs5uinb96nsQUE/NkAjJd9BcYoIysIlyWR0ixrRB6RA0Ls5XsSz30
ITG7jFiD66597gA86thKmdk8a+oRZZZp78wjruAar0HsXUQBxdZeH0iOHN7gV1E93f/2BPqcBaAZ
01Jp/It2sKO627htUYi+ERo6Pl4h7VSIMubm/cb01jC6DieKBud54Om6lIPPb3vuqVjpzdUT2uKY
0OTDY4ZlMjabniSE7PIabDQ9B1WIPfwWKs5tIEiAElbch9DYRoc/817UEKXlgyV9qMk73xOHMp+s
pocD3+dSS6/1VU+BsGo3zQMgec7kMXkk4gmGaPoLhOTBOfnJR20wIF1gf1y8Xfsq02mTNi/asrnZ
TS1327vQdD05YyyLHyjHxu9IRyf4F4nkZ9Yn/pXg9pFP0HtOcAAOfoAYhg2HIJBBZSumtVrh/3oo
vzrH+7M6LdH6+kYAq3SOWw1SZypj4OnW2AEKcgeNZekdbpHnMaMPrxzo7eKjKovH9gGo2LuZj1QL
Oko6UKAthO+8Qpm/Uiy3j9TmCHcqriP6kMV7TVYPgbDwOfbBAmVjiTNbB6x4bgBZbxlq8yoMKBEa
mEhlpYjl4C4AgcKgrUcaLeY8v6Hh1OiDzK5PqpqmO0pPrPNj8fehqnTUoShuDOOPcIi1sKUhH1yv
kLW/GMO28w73y7bwgycBy646u7r471zHepda37qkymnZMEPL56IHvZgb3/ADaAh6hvdsHURgr7uU
UcGnteyxo/6Es8m0DHKo0eM2tMyth84OUE3hcTGwVnsj24eIcB1Mr31KtN7jwQL66141uCv/W8m7
pKrDUPFCcMICBbLQcTRCWFClaPPgcNIFgTWglYduojGRGb33iDojW+9xH6rNqYwOfj324n/2ZfjZ
zqzYfD7oATsMamSKf+uy8r1oNFJGgHu63dflupItAKcO8FBu1fJ0X83GvH7pgEnkuFHBMRMN9DFX
y03tGbU40NCLqcLayQ10825OQP4HITvVzwW0PuZ8mIRDRnmsba5ulWZHme9Dn9Luh5BoKQn99wqc
Rqis9mhZ8LWadGnjJV05WEWhTulw8B0xviZYoP647zAGyvP9CE80M66Jf5Kv4fLeu6F89405TjiS
7cYaRaxRRT3wslBwYgjm3I22qi9UnAbC84XFhH++6qnoLwHsNfrMDPHpx0wM7rBRk2UFtr09rWr+
TkkXj9RECxjUYlJVRoaR9zcZkZN9nVu1lwgxYIsHDyuiEaDv6sIVxIhAXqJ4V2RNxPP9blIkRJJs
R1l3wtEV/1oxyfK7Sd05S1iE/7UHpsllFdLOGxuaRrCAkAkMo9d+3I5CEkQL9uBnigFDMwjESZOI
mB9TVcjVC6c3JXp639Z22FHBMB1WO/TDSkNI+P4TFBtrrLS1MK/gyxZ7b12MQFzs+Sr4+9CAN3oS
ObIPSX+1qSHSvrGkEpJxzLvLAvyYZ4HajkvUtdX7cBmxx5yzMrR6I3Cxfy8ntGLJVHHGTbERfg5S
D7/idmZeauiSFotI5RwERlgH+qcNCF27nGkbO2EOkoMXpVMxtctUhQm3GoRh9gkRS3USCtjP59J7
EYmSLWFZ436E2SxRCn2Q2RdcqW8uO7TJIU63Eu5PLeQSa1BVW/9J2QpjNI9VqSuzbANnJc0y0yGs
AqJEtNfwvUr1uX5G7lDaQK0y+Nf7+NtRIRySWsavLaz2qh9pQ66H5W57mxem310fs/3PtGn6fhve
Xotu+RFQCpycq636hPUU4/wEZYDidcbhM4byhJMJPZT8bFWTJhGMC/lH3cD9K8JY3fPvKDHatF8S
cc5GjlzdsJjm+fHtpIIXwjoVsEUHgINMJ0PHjLnJbqdC49aRNl4xVscNrghAKLUwuzBoVmee77tS
1EVFBLi/OpZByltEuGAF8U9SWGdSPbd7xB0o64KOQGt9Ma4xe/S77FrdIj4km8Zm5wgCFEmc9Ki/
OAri5rPbJ7JilsQLhhIJAoYKJ8R5xbKj35fNrYSqfcfhetnlY1s1sy+vqAqwSkhcXIufjVihN1HR
gKR3W82h+wCjRGH8Px5hcFT0TrQGvWSNU3RbHuqYRat9Cg72U0cyMFmoyrET9VcyAT2JNNSOTTjz
MAzQW6w/VJZD13fHNY9roujrEM35ZFtkuU8Xa7beDSlEVm0JHofV4X+RqedJ8oHQRoTRGrHOs+33
AHA6knO8SRlQ8GX7C9a18NxCyyhvYtdPoIzOKacKVai2x0E1H60tsNH5Bd0/8WkSxfjj5tgFGlwh
VxADKgc2iWvETnLWBqGwFW9VojOjPFdSQMAUlfTqd/uyVL4txGvPM2UUkDU8ukwneiWR524atEIE
3mZYk7LFH5L91lUwAlCArerqCuftXWlfnbQ3us9/0xUmQfaT4gFZs9K/mm1CbKbpHA4J6wcbyXSO
3UzgTfFeA58K09Wch0AbFhAm/fr+9cFhAdFae0g4E31u0v+PbYCQTwkOROP2faOROYtcCtxzvyhw
ghGv/oEHxdv0PePGCfzbKreydyD4Gcq8FiivXvoYzpYfdhdbOm5JaC0m/SKuN5WprJluyLax/2Qh
5oizQP+P+VpJkOrI2/45yAOlBwbjhONiqkJBfGGtX1bJpHqRT74GYXs4jPVmebWu4UuYYtHX7WY5
5OILDJqH06xRlxssUs+7dpHo+qFX3KGDn91nkBoSbjZxUyhoEzc8xyCpFRrwtSRdZv8cpf0OtiMT
ktL0XCLPgTt6WAMUFAFohz/a1SMXc8yqZyUzPJz8ydktYJnjB8p8dpzj3QhZzjivrrMaT5VRvv1S
wNvp2nlhKueOgjFwBUDKAMf9nxKFVJEH1dkkQN859v0X0bKVnSQGOYHX0D7IdzuRi+1HKlJ2yJKU
/YOq1GRbxX782OPqT0hj5bktPLiZHJcFd7m2YGtPS7lLIZp4wFbHAxh7BhsrrvdyqkRFnjSLsQFS
xsYQJ5KC3089abxrTdqbC/LIWrVTwNd+0Rnl9SmE6QRVeYIECyxXShsgivkj+7rVbhzooyICD75n
8GrhAMnmbD2oY2jPen98NkfjcJQKuDZcM2SEldAx3PyvQ6teoia2qJbWqpmCYIdDrnzr3VR+CMvm
k72suDZUss7RuhSwzdOIyfD0rmaVRd4uddPlnhRoJapIT24yXHT/oPRXYAGSc9n7fQTFvTfXTVHk
UJfoIkkSzWvRBU6WNCobuUGSU46HkbmzsIsqTAjW9tk/rEGbIxzpNJi7W+QHUNJyb4BR5vuMURDs
YpiZwhpvdF+WwqIe0dz2u7hb/3zabaEmY0cG98ittVc5bUCJVosvD1iTzhi6PZYZBXzyJS0zaRJC
KcxQDKRzEk8SP+lxhsk59xkkmuqzTL0XdoHQq5CRLXdbjFU6zDJcy+siPbiw13Rs7eYY3yfZA08S
QzbdNJKzkq3BRxztRtPzVbQwA8cT93cT16cz8Rh/gf1LvrIcZ/mbEG2KCkzuZkVLknP8wPeFIglP
UCkJn4Ffl6mcLm5DV4XBadTNaqLV/f2y605tKZlnQZtWH4NXBj5jOx76HTlqe30bGqReAk3f1U8O
40yKSgJB4Rka0pWr0gGt8QKiJ0jlM86VKS609uFXY4E331eZHqNQkpZukgOoz9cKYhw0FhRscqT1
84AvmCF8HB9XyDmuVFOldcl7CvYmU9pcIT53laELcvoVF8mKi6YkXdfrmgG6xvboK5qV34dVit2w
7sELR0gt03fvpN3em0R85yGJhg4T9tXOM/5DNf32pErkrQRS1nlpItCQO/N1CkMmxy6ZeCKFRf/l
h26+0DKnOQ2wyFoIwpzsg7V7so3nWahOYcd3nHmx3rDgkehQcpPQIhS4jOGTtxUTJA1yVZWvszsx
og9NPkQwzrreV87WWSkvwi2Wf2/7v+TGpox66OYC6Eb1YSqEmewn1PPna/vP2ynoneoFnsZR6gAl
ZubP5Wdiwj4usVgnj1BCfvH9KGXt7oZOeaGgOjT1W7yJI8fOLjYebveR0yinz3XP4L5ZVPEcjxtV
aO+kQPea66CgQMCYCn1jkR1CAs2qc4cjOg6yLUBk4BCZBgwo5i+WfEe+nhPyY1KyjMY7+9Hsi7Xc
XIXwdzVXG1nkwyadmS1ta6OHAhJHtkXr3yEoWaPyjWrhENnPfhBQlGFyoA6LY69DtVZUq9iVHCHO
HWsH1qh+x4+MKcH1sJahsrsTrGkA/ZLmQB2bPFFb4QFVlbCDt4C+dgPLKVvFGxz5HnEMM4w8NNw2
f3FxvXwD0RKxbhgDVliR6nHtuDO6NyvNH/dz8gqLr0WjcmZ7gfwQOQpMDNowDqs9xLuJ2lrN6555
pSZRlNeMk/Rnfd0NPgPN3cL7sBabK08t7dDmgSX+UimD8kHHJP1sCN1PBdVZVI+Rftuv5t8GG9Pr
5lmBUewGAzb0/eCdDyHhcGSons1eqsGWR5sLzeJocCiSIfH+QARbn24GFqP1BdVvySRrYIewRj7S
RzwOUVtUxJkvall9otA13t/xdl1oPmaN24i439t2leWq8HYGihmqfmmfGwKvo3imqqCFqDSdZOpT
H2FuOJdckebcFaMNWtr0+ACN+/wuk3rpiXOamekka9mVR8jSDzwFF+jeCLTTjU7fTn6tO5pya22m
KZRQRGKfAnLSdQtzCfMNS0N4yOiHE97VcKBSO6VwiyDFcO2+86I9Qz545SnzO476A66paemE2MH8
m6u7H2sjB1qv7W+X9+0kEBRDKXNdhgI7MMzm1Dv/nv+7sBCuhjSui9nR2Scy79Ct3EBl9oV27nIn
R85kD0mboYQa91dcGHP1Zid4xLng+9M++bg9xyzY/EaOaD5r8mwbEzcooc9JyUgnwX+z1IBMCqYg
ZlMGHShZyUVeRL75Oo8WW8CqTrmZTVlsu4Dye73IguU1MEoFvhffRw8AbdCjEGOM7jN1jirFNt6E
fDsAGWa/AY9rYFOooHTc0pG0ZtBwcTnQRclKenihHrXMhFt6GqL5wPpQyubyKJbE2CrSQ8p8SDFw
cdabLyRXG/1ZLGNS9YcsgC16WruSGwc9xu2fR8g09uwOAaPlOVarHj4MLNqTOlQSQKXEMmsd4Mc+
Yc0lfXybmF1WRh1klvQhzXkWqGbdJgajsCOuaCBd0zhJ8etHq4psDoQbI9tompEr2kzwpLWgqbyq
qD7UOf+EtsvKaJm+94gv/avWaDLQyb3lgcfWNbK+ZOFzABU5PLuY+5rF0bf9O6zk3qIQKmmDW+lE
73vhSG5wiMlv0NA23boaiMS9oCHTmxiKV8EnihUnHsW2JsBnNfgAFMCCgsAxG+7xG+ae21mI0F31
MQ1kJE+3nniuEiTMA3bLTd2CASRNun7bJshv6CRgSnaynB7bqefEEXy5mLwDRtQtSaK3RGN0p4x1
ggWHy83NBFqRGJB/N97NIq8OLqb/72yUTUTmy1I3NaxL55K6uw8a+8b7X4KeKjjPwhjS+kORzQIw
TcicXLYWJOowXlIJri0MixbGKL2Jq9vAG5zn75rzZZIQYZvyRWS7903ySfPd0I524ltVBdVMGvJh
7SQLrgFEkf8KamvrJXrTLZHxRUEeBnUiUDYq1GZAsgbEawOAZ9VZwN+wj9tc8PIq7C64XVqkZb88
0GLXsmzqrO99XXfislZISk9Llj0wigcjK4xOchQXH/gZaVSmDD1GO8EqnJhbeEvRU4g+x/tLOJyW
iXac9xGccGeWGgcUhzk0AYXgratFm/pdFm+L7w7aVbq7sLuCLB7duDiA41oLeTCO5qySWitUlApY
32eWM/8Rg7LLBFDBGrRxgFwUTgFohu+88UXq1OhS7qLejl4AQsA0p0YFbTHpNOV1WrM9Jp5tDzC/
P6jo3uJUAvSXEOMZGiqymWSr/ufw/4ZkAwkmKKQNKOLbKelaBoxWZFlEBK83g9Jw0jd0UExiUUK9
WjMFyD5QoqyTIJvi3awkhOiI8l36QYiBYsGB9735LgqsTu3zrEjDqKl4leMEyoSJhiJyOwjV2kxr
WoAIXizniZ5/fixYq8doCNSr/4zBZyfoe6Xh+n9RZA2DvrT8tBKF5sX8bcGrII27PSifxO3UuaWx
kQqfLguEyyw6fEjjExK/aJxNpWlG90OJhzq0oOXF3RQ95FQEZ3Q2+8nYBduduvBdrhZVemYPyyPH
AQyhTtwElw2QTts238Lz1W6HjA4E2gq9UmKMtwJZHcvEtyCTvnAcQNd4OJ5Oc0xEMH8/4gopS9Ab
tdt1odOhA9MOjVH7OcISnsCEQHsBwcXVl0mvEzlfFI9icf8leOtdmkBj/AUBp+CYy0cmzJKwz1GV
asUmLfZTVYJhIgP0Y1vWEVTf7GaeFIi7Crsai5Ud6Fd70odPRY8cOKx6aLIWvNdeMS6oS+FHVtVi
0MivPM8X+AL9pJMnZi5ncRl18/trHiEpeerlp+m0imnIsK5NuTm1O7eFSJxx5RKaWiEK06qriVJI
Dz+1blKk2VFulxW/NtuCq5PscMRRUfB75PU5I6rlQJH5aPOJUP3hbzgRY9DX3Y9BjhT7kgjEefW/
wS24U0LIOPXhnVOpqqk5ZZBBohX1TxEEZwmUVp8XRHYaJ7IHxSSG2YLz8bSpaTXTVck2M4NUCC1M
OaW3lf6q+uTBehdWZv0UiPQfs60aDu0KrLVtOJHexOnkEuw27UOsFECAztBw7F/fjbxII5WBZLJi
gR7j8oHcFdQKddCB8yXwHgQp82Oj/j9ox2cGfE0Gz3nec7ukuks7PUED/vVSCFAGca8mYu+AcRz2
YLe4mXgpW6asDSEjs+KWzVbXAPYQhw7MizQajpd+53LrOsH7HmHFN8YOQNjJNX0maMTEnvKBsnPK
ltrGSjpO6UE6tHDSQKX5zhHpjMXc3hVS1U+HgcG1b2ZDeDiHraopEM6SgQDbFJnPERxuDviFbp4t
4EW06xC8IMNtSXsLFu86ML/uoZ8PzpvB6ugCKV6VVu6Zs+M/qDhczYkLqzcxi63Uz/clRAnQBR+8
PzCksquUrRHNyFoOqg6A5ut1UISA6o3p+EaQMzlHBTZmG5xXeaTLSlEjZ2/0eLjxIbQ5rHct6d+2
7b6gbcPexC8HkqRYq3U5+Zl48ORXqMWeQmm/zL4j6kakigNeq4VpeHqlRCdMIYcdmTZG2np77yag
ZFsk+p74tsgP0G10bCmNf9JOCZB4udYZZn81WebtnwQA0ZwIJwONdkRL8zaClAe6+LdJ873vXCmv
Aprgjv00pVu7gQJsyxICQQaLrvZ4XwYwUo4c8N5P6qKtwYgy6xVI3xAYes/SolGFC6lflQ84RhV3
/4reFRfD0SGQb+LEMLw9v7uHAQH8FiUVairarEuymWkcmYlJTcAMD65fITBgT/OyA42U0ySDddfI
RJF0Pl+Rhd2RlgBiIephhVwStz5s/lb7QWyUSoud48hyLnmApVreR3ZWi3gGqTNQvHmYrRKe8rIF
vA5WlTOj+5SnLhQqob8Tp8MAFtNGfllKSYswDrrai4jXcDMMVVM2AkWNMP6QtW+DynFZoN7kR2DS
huBdEp6/VfQwjHfV2rh2psDKIIm1r1xL2mCWQeZjjxBeGGvUD8UxDVBoVsdTZhfT1JLcWkX1MQTd
H+omp+UhmjtbjVAjXYaDa44UkwkB8aYQeGo3LbSyRl2KhhAMyBzRts1dN72zYTDEHBycMurAX3LQ
VNoGd1eLdzyhnyo2a3AgHRoTgOVxvWVjqyd92f3yBcyMBnYTwHX9txVfDrkiUbr1EuM6PgxSMzp7
dnW7z1c5VTmSbEmft/DPbTio3Fd1fTrO4q6VrXOgFapueXHgOyznZ2G+RfqeiftjF+bBeVVq92ec
J1C6kVi7K6oLOxuQbt6lSgiwKNcAbU8tTfzZJjVuioAjBgsiMByHyjIVk4wsVyIhVgFwlXlxrA/n
Gp5eC5z8N/urvIxjtuZmddQXtObpEEjnjlliZ4MOAPc9wuUhEkQUPucpeJz/Z9JfNCOrzbaX/K3q
JghG0WCwL3zeE4kc2xf3CTVdVll39bzpvy2yW3Vdwyj/9+uIBsa/JfvFMSq5zwt0ymX9v99x8Vlt
iKj3Ww9twEmdcxjMTrmvD2XYpUyT+2K/6zFMpBS7ZRclQR7VOK1ySWRf1jRI8pcN2/hCXX1nI7v9
PbDkPyl5AbQWtaT9YdYtv8E/uqOwqIHxeR7XaWeScPvvSuX3S04N4mbIHM2E1jaYDcBmS7AJxZQD
Mjv3JDK7KscIDCrWEzvKBSTq7EnbZpuQflJiIFgZFu2gmuje8qS4+0DmBDetJ/0Px+y+4JpC19so
MesI7BBT4HJhJlXRnA7zu0e6qQn1i5Ve/FTaMYh//v/JRmxU/bbjQDZLFNzH+WhoUdYgN8ZS3w/U
JOrey3iCDCkot8Sv+ex776VC70jFKEScZ5+RJHkSy8SCYpqfNyRW08qXD3RY6e/16IUf8JK8fn/i
flPO8mNGuk2EICsqj9vy9JxsE0tXbMv/Lw5Wklp5lxlxB2Vw7bmsErjS51xe9PnuNK/1R/FMPsd8
UUs+TXcEuzRRSHozWaomktXu+bc0wBzONkOknrqvnE1xqkSOB8uQ3Rhx5Cjz9hlkkHCK1dCBKVNi
9THMdCw3gaxtiZMOszFOsFDNOSHcAkB60bsPQ1+e4KY912862iAhrU3h0xfV/73M3hoaOagWiuZe
oMedYO9BOEBma8G6abNdJn19WuAURu0p0Cnz3ua1OnYIAS7nJupKypWRZLe5pk8o4YQHajjNWygl
0fp38cvpMRkUyjcPsSj94FoQ3e3S+bVWvaeYhoqkCbavq8RJLXqSektwJq5icWqsxq3pnJ40tM8J
AeDBx3NGxmJTFMd9wQHUdu+/Lf9AsB5LL8GD+6AxwG1NjntyzaRwtlfPQeRcP/jcLwmeTWU+Pwc4
tjiZ0TEkv52dYvpahrGrCITII/UaY7M7VDpuW1+1QnMc7voaMbm1t/DPP/a5Qwvl0LbTE14XzrY3
hQWKehtM7yasXVmJtaS/zafy66uZmtMuYiMt10RoRyfxrBX6YOKQWhqg7EIuWMGWbAVh7kVopD6c
67FqCZEPl045dS1NepyE5JAvJsjj1rTUq0Yy1pSVnzcO8EyllFb6hB0z0js+tOoge7Y687RTnNVz
VMjnrC53jCapU8E5/zlmmLnkNkSZYn3lFu30uEntolxGpOOl6DUp7/QuxRK2ayPNKeegY2mxlaPj
J6Mz8+P4avXmbRRfKlgeJOuBpxX9a4JDsfU54sVJ213oBNi017M+DMCcFN87BuBdkcYfUefcFXiS
eTrWlTmHM9bkEzmXbwRIEV/QwN5njLbyPTXrr+7kb4a6bwEn72pLZ3W/+sduYXpktXxZ4Hlqrncc
VrJ/GV+0HvVvJ4bTvuFO/eTyTY7QhpuI/Fz0dYsnpD/BpN+6OR4ugqYrx/JMxEORQX32wDFJuHPj
3OFOMHwNmnLNyn3oePlXxD4JrOXs+n39+rmgO0hNXFr+/mRBGJYKyroD3H6bbN7qLK8cD774uDhu
W+Vr0Aqxn+8g7blMwDQ7Ek0zkuwvNY6BRBsIjq8WwJ1xJ7Q+6mr2I3tU4vQRREgcLJw0x/rgLXjW
w9FuQy3uRytVlDYON/aXqY0bYaL1+T/W1hIevELMsas00+9XtNocLxi3a4IW2D4o/L+893iOe0F0
wiJ77yuLWczOtm3wF9tReSAOlyrQivZi8LVmt3XWY/sFIEmnCRdAv5oJIP+vP4n32sKrGxC1udSn
SelxhVbqtyYfRBso5D96BTMeMM4lE2QnFum65YLq1tNOBuolDgrSLFg6ppVud2Z6uXGIzEohgOJt
pXdf/HxWCRD+6HyWu6CTVSQcABLqLNmr0yIZ/OGQ/ECcnwr7K/AWEs/PFCVH8zjHmv+LdtFxG4hr
li0guiWcpRc9HhUpb8O/GN9FoJpWNidEkATFgM0BSuT7xIj+ImPWpQIipi5xLz4Xj79fNr4oiKNC
PlhV+LSE/y/SCM+vVC2clCZfMNlVZyaPeLOxr1KvMlk9pGHdKjkS7VsHvRc2tuT8n8dugSUx+HSa
tmr3vBijTZugq27Bb9XaT3jV1XQXFvBXgNtzePOrcCfVtoVNx8si41RwHkSelc7uvvzs6QIYnetB
+kbU06q2b/rtCzHUyMqQDA2rCFvK76o0AvVQ2E7q+i/uMKoUU06umVY3zMjCNvkyZqZnBef5rhh6
qiLdGh2NRjY1V51OP3tMW+n6Dckslcnj8q4x/e/v/K/DJFYd8cQh8qst+IBGEuMZlDaHkTjYq6MF
HRnByeSttZFBSGoTVAfxRyRywk7h1+5S/lHwTlfmzq6C3dTBVHB5PMQ1wR1P4uOnGt4lqgHWslB/
wA6pMPJGUzKjtCm0eMMAladeKmZ1V+zeQHYd2lhKdWTc5zQeqc1DizpZGDszLgkkqYtqMaFIYgbb
jVmEj7jaUZF4R6ykNp33FQMESgTiq9Uh5JgKkXVeaQJA/QWJkstLpdPdZ87PVOMthuOujaw9f8t9
Ip7pHp3xRP+WJaMfxB6yjX1DKy4LaJhwaERB85T4UnExAGCMsrL9ZYPHiDOJDLn5kJLIU44ncLl3
pWXsJ7+bx6YvpDmxeGhNeazcs6rcYQA/eKO6H1xeo4yX3Z8mOdPebxjdqyzxf60XrXDIBTma8B91
kn1zK2LRV6bpQxdnlxSukMgnm0+6z9jSvzUbj5jr/iUvzNaqFCcemlNaDqkw92PJiVZy7/70QBTk
UA+lm5L01H44jJaCp+e532hAX19J3Hz/dqff/dEMXvOeIkccwftSL7aF4jXjKy34ikLcAFJEuAi5
h1jsZJW1YH3TfO0sk6+pJ9Wl6PcIw1AaI1GBHiRWbK5i72HqtE/M8oyQOyJhLqHPt7Guah6TpOgd
winOqwnntA4yOuentrVot+6AWfOKxzjuZOQQl4HGYadqH/XI2AgM7sOlSyfPg6jdmnJswRriEoQD
Mwlr+zTaBGdGu19mNq+7vu4R5KlbeVhgnNxQ9zYW9fkhanIdjP65K+UGxt76q3UDtBXYc1O2EqST
tlXEgQvInwu0zcpNSiTB+Wwif6qcmjwfO6JBRHY3gy3QNDZ5ErUhOnkwsWoPYsD7NYPaMb8eeZz3
WeZYJmGodSY2V2bahoQh+UYNxxfwH0M5Itdf7AX3n4OLlxeDBRJmfnCSGYZfdSaKluZ5ZvY/TpVr
RfEeAHr9z1HdlBsECDCAW9XryUvvlZSov0GQafJFadQjHvh2r3Yw0xtD3kIGoULtImaLuVulnTHJ
qDNgk+ZoCFy+mNEHrG646tHZFCi9SpifYwqC56qhoZFjnP8VfUEh4voZPXv6fLKx71J6PfbY3YPZ
OuusXMo1voaPdEbFMx9lKdsX62mSNwkDhrP0U9ugaPQ1mg4YhD5DXexz4vSXja5t0Mk4OhfcD7W3
UmtgZp7KSalz0dN06sSZQZlL1XYQicrOjyXoZk+AI58y7Ld8hmiaAJCOjhpie3FvOerFSfW6CzeJ
oVX0aOlqnx52Cfi1ElER3/Qg3ZdD3mHOdD5kcNYUUafg6M485zgXM1sAnEB8qF52YxFj/GWsdryY
RQ2SBmoGFYT5+esEtQteUQG7NMZgohUVr1rK5t4REis6CvobEmXHttx/Q8qpDGbVV3NcQCuQsU9s
IHYNY1czgQ5f9cSEr8tlatUyKUzrcCm+jd+Sp953BKEc8qcmFv/YuZNWibFo745XwRg6PBge0/1K
BBdeoZtEGbKGJExpfYJM1+olyKnLmZCn9Xie+Iu8HR17nABJTI+ytLl6SLCABjh2NJyO110khsio
xKS7busUHKetT960l1XktkKEFuNWHOGe8ojKh89DvkV/NhwiaN4KCYzhM23DySO+COipifNBHlu1
E4G3+TsXDfx7mbUPjAGF7wEGHY6CDve/zmn31rT9BKeoCOyxlsxwNTeAjynGjJk7jBl3/4ZL9Wb0
2weXqw7FKkXJlv6thX+t5ddwY7DsnnATxNNP9QGosDcPET4eo43Eex++LdfO61nmKtX1nlrNEvAE
X8PEFHAqgI32LQKsuk+Hv7bBfxypfCm+mejmm1VQ1KHEqqjE3oNRynaNHqfAz0fK/r2GcFdeJBzx
PDWh+pbXsDueafD7wS52Rqh/xNaRchVqlIpgU6/Wxeas6FyQGEFjXj4bByaDJUa3TvQqjPEeolu+
KRh09y0UUQ8PtVEQ5KCR2fYwF/2mmWJTe7GTVh+8U+erH/YcsmypslH2HysIuTuRGkiwJlQ+BY9C
fOK9j+QsPyklGfCvn8Ttdo8CuVrtEZpOdQ26ZegEEuXrCo65GUeUqeD73Hl+I0rNXD2BpEBetToD
Sc8pj5gvbQxUyME1SWVRLFslXUxJfX7aAboScmKcEkU3E1fNZ24RgYU5caNKp0LjL6GgpzXOqZ6p
f6BfVV/u4tgb8KIme3lKVYk75aNKORVUEpTvXK18Ol3IrIwJE86Fk7B0za5HpgpO2SisRcXq5ted
knoGrqdaO10VdrQqt/O2m4RXvRCUtlWt+kGuPOxoYqJDNPgbjvOaHBQA7qAcL6yUSqDPKMx2EmAh
f3LONL5SPI5uJpfDNa6HN3mMeGb+/N5Jry0O9GLpaHh8pbIwKUPmnxyQAsVS7VWuQ430xizh1+mO
H1bywd3GTOyYz9fKg4OM2p/zzf30eSCFCRyLgQBXump458AMQnTERO8x78ImD7zBAZagEBVsxnoq
p0ApqE1UijUGK6SrsXjgCLjMoOEV2+i+ZTgKRn92YcZY3MFLd6BqKnsGIsduahfklhrmKMRHFV8D
kXKcMgHkjE1slwSAFJ/W6UWzCt58kGOylGHDxVedvamuUMNAavQD46pp0w/nhDrfPqCAmhreVORt
FEfLywTWlX4+AeVMFxMikjbMqROmXjSF2EmoYXVIUk3Gm52XBGBVJGWEKdsfmJbpsUpTKXC6YY1X
xoW4TzImux/Xx2jpIl+ibucNg1n2v1T8n14gMLShquPz160e77ldtBUflI4JeYj5BNwGrnkMXr/I
usv0+lbwHOUfHpNwWDvvpcBQAPW3fHzccYHR5Ovwwzwd0QgAU/v7+vjnSkroURzGDdTDFFxrl1+M
VxbbNqNTSPeY/ZCtOfD6qomGgzdQWtdopRgB9moTX4rrUp391qCMkb0LxL9LaJY1I0SXIhVXrkW/
SJ61pK4011aDquGWRGLewp5ddjBk7SwhWRUfbWyVXl2/V1ai9chCjWfDxVtj9vd5OEoo6YpLlN0Q
eeUH9CPWiVboycbtzhDjXFh47K2FG6/tQgGUZPjcJLgFfkUcMhQEwVtbYnm5BJcoBFZxeyNC/z16
g1d2Eo9P6DUtkvab5h12ZmjTqOUqQ2QMGuzEnCqkpFUE9MBzJE1Jg+hJdGvLOBJ8ZXJxBGnmp0rt
rJDZD3nJw+37IOqKlw1Ofx/4J+7fat0TVVUpC8RT0tuEjs/WQD2MZ9qr/46+e1pZNkxAoatMVWxw
6NrfTnTjD3Bqbp4pgBodXz+ehLRTaz1rZ/wPeM51onTDDozPU6JVoXQwVwYkGTqctTXIkCOWFYrJ
50aDYWgSVqssLEULN2PPoTSuKLU8C51Af1iBOXVQe7CW1UdxqOPHvQ3ZVTQoSC0dBgw9Z+rzMeRY
sDVvg6SKPoT58qm43yIwyHAg5VYwmqDsJULbvi8tmM9NU0QeQ4q7EuGhL05xjUG3fV5RzdxsHnHo
NoK1zf2+TUsdhMD0ndg0+kcj7YRABUfAY4/y4XSORNDqkgsNLxmly7RykxKVOd2Cv9dJZb66Iel7
TGK/0FxYeeO+hmbgmkPFLusKHHhe/Ys8cmoFKw5Ytx4didwqUMgBE5J5Ggp9PUaQWFPjPkIY0rTq
uC8D7b0cb9WeQePYXZLWPoncM4BxnzQlTAmQnmwQ4X3rwaMLIszgrxVhraaKcChByewKZMPzw51Y
hmb28Zw8mdy3XEnKByHavaTEia5LOXz1ztzWqvROtercNw7cwIu3wT8iYDAd0OG9uUv2Vd8bI1E3
Q287vkXbiBpUy52bRbzDd6pYWx8dCepTjg+dHmmBzRGSwTHAsAItUTtnQeWRG4IXB7VmE2x8NDtH
2xcQvRFX9yPtpqbOcX0aM1IrsrkDU2t+d6ljW7mjaBm1NmmgI0yy33QNyWfd5oojaBvZAfUljn6n
0S4zsipoP9tabHfO9RPr1iuakJG6dAgW7g+v0ROlYCQd0rpqwQ48qdtXoRiAbB4FXUoa+Eu9JepJ
w241sa2vPt7Iy1OLZgRs0nepC967kZj+KLV4AxEf+zL/EFvjqIeXaI42JsWLfhZndBwusyIt6Jnh
QgqQ7ere9qhu3/N2bgZ6odO7pH2fGu31UlMvQz4gJkR3+viU4+94qOp7ZvVpyhgTlfofXez7YJf1
KoBqri7FuW6qSsGjuqM5guCTvugZLShWGFEqW3kvPJZVfTCkG/YXsdn1Niv/9ZguNCx8N6Wd2xaY
2GZNbzlsaoxfUd/uhmcAwbxHZk+3swv2JUaIpDnwKAm+3fzOHSKBOxwZIgD6a55q8rurrTkagsx2
VxaRVc62j1Rhm4nszwFYWvKWfjn0lnG1pDmgpnQTN/8rfWWRRcq7ZZ7bQH+DG3Dysgz+UuLr4pjN
ULmK/slI6fPcsepylt9RrPak9nPaSgsCH07hHrUBU1bQ+dzhZap8m1nEi1TzrSk63rraTwi8mxVp
Q+ziC5jARmQzXnojMxnv0MvUqD9lwN+fo6/J71So+hRlPIMd1mB66e3Y4gB1IpAgTLJz+2ld0ZXA
MfeymFBVW1obj3rN4m0waRpdq9MSKcW6qA+57045rCrsnD+R/DmWoiy5LsFsBeE3iu7JAPO6tAg4
7SpvGC34WHk3eMFP7rqStQXSWWCDqgHl5FaM/qUndDZ/P0caGKAavjgCYyu/yBlKE+Aoku9RTqcW
8IONz3nx89gPNlKapnhG98XhngdGSu1I9yLb+Dn4GHBbjJdo/W2b2LBwjixYVLGfBMCFxWiJvXLV
ylQkb4SqeULdnPwOgJ9FoIEqFugR36PrRGq7GlU79i6DmHhvEtxFW7Sq/YV1++6ESsHe6uVTt1vX
l3KgyAg5zEnTqvhGPfIPATwQQr/3shPy6gKva/I+VqqOi90Zu4L/rFuMOfUzmmwEAkPgyxlzZxnS
iQJ58l/lBDtz0e1G3J4LenBHKkeO1d6GvXzUqfzUWVLmwb1lSsqX7kF4iMGmgIjt330c4Du1lcGU
PGGpqHidkIBdVPYOt+vM2WYeGtTIo0f8qOSK+O3lOb8SDr/l9wQN1k2TTDqpnnNuSFrsXOv72kwQ
KbBpMCI9OHcgnhm5yzk34Y4iF0RpG9/m//i2wuu8BA4LinTy1JAv5mrAm8aYrDl2XxJO07eGZQWt
cejuh7oNQXyL5BX4flsoAW7LQAiz9ldDZwi47C4zClMiEuPKkUeOSwvIbDq53u3y1j5xhjoJ5v2q
hG3qzfMUWpzOWvRMK8WutnKA2XeYTZlas/WcextIVGQzWnqeIli2umEqUehoBP954+bkWEdqLAq7
OnYy+0gQYcJltUQA9FQHwzXe9QmE7SocYUUGLzGTwtsheL7Cnc/lrc3wccF7Jd1FD+jrLg7smO2r
2XjqQAWDFSybgwchOos4vkZN4dVJzwJJ/+xzVkYd7UmQd+2pH6bfWjc9GWjrujJqH2tQMv3EsJi5
KafVf0mggWt2zV5ZiUKJiGFJMbR8si70SpsRy3rl1S012bUvq8hqUPi+0rEp0wqwal8LkUUwbUyT
0DsCBCMpVg524Te6Maypt1M5Qz7qrpolcCMTLSzWsxB681RrfOcz5WyM7u/0Q/y2cCCGylsC9R4V
+ff0vOGGSfj/UZwrbCx68M24MKFDHQr8/1YxuKhlVY1UuikAGBUIXCOnYuU2sq4x38Bj934t+tyX
DmosAHByb/KYGXFrlWlewh92HwcKzjraRlBChte6J5JaLgl9YE1CrpQcu4Os246EURxrT9cmDGkv
hrxFcgzJ8EfGjMXNaKdvOR0+9P5gVO+RBw6j51CGpAphh2VW2JxBOu8dK8vOqGLBXjkYc9LHDPEj
5IgHM1PgYZFoOnqnB+Khv8rhyYERAThQqGxQjXhMPABia2rFPOKvB/8J0OMq37oa6U0eLx1yGWlH
rfGk83rQD5Hyrmj2zMJl7An9wp10o6TXfN5dO+DmlE6BA9qMF0lQPoIWO3XW0vOjdsK2dNbY1bQH
5R+efL+DzjefHgNavqXatmvRzUb2W+SL2jFhT18IFDsPHqy+ThYJgLr47yTp1Nau8AJaRFzs8eB+
u36pRiCpxHxXfLyGid2956L7Gp8tJVvYOGx00rapOqTAhP/ZgrOXM5+0CuJxRuCvqu/K02awHtO4
y81qi4zMIe5Wi42OAP/7KkCy6c1RQyW3Vvi8d+XKtI+RoZg1VtVscxFWXkt7wn0uJjYQLUHujome
8dXWDzjlDxXk2FIk71N+CeJCJK7yn3M4tsjEddGtM/e4MGU60lFXpRfbCb89ZrhYzQgOMPqGiR0I
371GqVBEeoh9fW4zNZPCxs36iJWW1tfuemJtL8UJGBDgCGk9nm5h6LKfuNLeTkhSQaL1nwDAwBlZ
nRwJmrfabn/vckikvDbZdQ5wwWjx5JK8fOGigu8lknz9SmVqoxR8p6MOLdPGP8uA2COvV2iFjloJ
MQsGupRNeQxAIO6zy4J/diOmPb6XEOOSoDnDc59aZlVQpK4j2Q8QM89VfMK/mlDr/sIisHx5VoTe
3YtnZm4M6YHlkvt51vKOj1kZZH8jrlbWmIEUtfbWwx+3+ZHRsvgcJiaIFO99DpQQvw11B3Rp7ekh
/4B+tA0GoV69Lqi+azDgj3DGeOL5+wSHblLbTqxtKykhN5kBjEn1U4UQ1TTsMWfeHBddOgBtjqwH
fkUkCwCDgLVP+MGQVANfTOe//cWFv/JmhKha4DuqPhDh7londvGSkM4x7EHZw4QO+AeY3W58RceU
CafDPZGmSFQXTQ7gvQdOvXroZDNcWqlDD5ytBaeGPQpech0GoGKNdYwP4+YGMSZYjNvSPdc7VrV2
5dyKDyv+ghV13FFakYJK/w6T7eRaZotsL7CK2NrdfK7TwDmrXfteZqIFzhIQ0x9NlaaHIxnr/17Q
URPmgebUElXv0JqBCgTOH8QD+5ljzFUmY9WTK5VtoDSzE9mpx872+qn7AiaKL7PT/Tw6TZwXsOuI
8KXK2S02bNsNTMkDy029f/EXnszYwOzGB7rV2lvevtpUblsbUGYPBcKs9wN9rd3ESfLxZ76tGRbd
2Tx8dMUJLfKF2o21ggvDVIgs9isYgwuUBC004ueHmKMeo34xhXiIaM+lhcMsMu+/W1cXuQw2iFKW
KqMk3sLp4HJdJCMQi/oHffL6lQpWMDP7K34mcAZdnhizLdtm9/Fm5f6Lc/ge4Jq76K5EEazzwQsd
NO9aP1RceipeGqvCVZLVEQ8VXBn4dDcmKajabdQP4AGmv3MjPl8ZsntntHYRbacQBpIjqfPk5iCa
BKOcl5G13jquRs2mL1z6ARpCUZheSn23DGBk96TlLmHXsdYlJ4anZxFSWwzPGMH/6uHXYe4qCGuk
FjMb6Sf2f8uc+dZzrXt4BwNWg8KJWocx7dN1T6ItuCB3DYIrTqpWg9vm7uXaasuoNBCLyuNAM2I+
Pjvy4/1YIfKKl86L5tP16PUxOcwetOnK/LbD3NqYYEx0p0/ZiYVWaqXM9NymEpFsTiweLynfxLZd
CnOOj1JchhGdq2c2ID4/eZytgtdGjND/cDjGhBCe0nHGJ6hyNXYWWmo7kg0y8EJ8uv+7SzGl360O
qCXL0LIvgRSFQln17Lj4X8lEeBQ7n5CqUAAg8MycuYFHpltkrwoeut+2JDhE3Own53Hjz/RxiNvG
UV4ppNaTWZkmEYBukYH1oq4RvW5img8JBJe1airn6kdQLC5Y85rnUI3e3IyXpX86cvvduX1n+ykD
0NRIt45AGUG2UjCr7VXbOkDp4g+e9Z6hcc89rqhQpmRhvmAxnDDSQ7nJgtdZX6voOgo68CMkuJ6H
GFHk+EeBl4XP3sBJDPKjQf7ApsNMGRtbwbVj3nzHtk/GTWgJl8Yy7+MeZ5NXLOVV56O/4x7UGD6n
xlQw0zwnAQle4Lwj9AG5XvXT3xPTlWg+pcPf9+z398cXh20owDUzxH1fiSFlpPrjAr08nLqK1hPU
DcfcXpQ1xAZWWAOR8PXap8O8RF2VRh91Y41hpjRbei0RSntRwxQAiTyPHHWEwVch4yOnD5y7sltT
TiNamYp3SNVKnRiULTmDRs/l0mWf13VdMGs71Ao9keqyGHhzYbL62iw3ezGzmZNxxcJ7HMOm8snc
FCSUQ7il3jQgkkMwGWUhFTwYQN/53cSrYpJnWd3FdDZrLFDZ4PmsMZ0K45f1defCKdJMBubfP0RO
TdGAvUt2mqx8Qv6ZNxgBY1OMhBtBx71aafmqWGdwcGaZfaoOR3C+4EhgByrpW3M3vbpWlbL/oaN3
Wv2kSw0hI2BsdG2i/QuFoh0DTO3baql3BVxru9CeVclFp7auOeM7vT7xvDvnbtBWcQV6w4+XktLp
7aDnb8LpuWkdD4kZRsIQtGz9xdFMilvLunVS+6Jvp1tVh3DIoGTkFhoJUeTnXnpUmRWNJ+oEC3xf
zQ6rGL81pdCPfzqC1657MbJrHtQSVWYBZTkr86uG7eU0qAyBwZh+LCjwidYAVk/B6e1SRAqBWHF5
zldIrOOGLkptB8xS3e6Pwx6G7P4+5Ee7RStzmxHuZHwOSxAq1/ADIY7kLG8hrCF3MZOClpjv+wAG
FuauyxDjgazeyquk1o7bb5cW9fRI/M3cbIqV0vYEKMLRMBuUvtudyGWNg82p5yw9AkK/ygB38ds6
m93QjAagitOxt+VeEioikcTAUCbHUipy1nnrnJEYI04E0DfG1rNJTGKA7chi+mGrm4ncQkep2aRC
5EVjVjf9DXEiKb8CJqdiZENJ5p19yA1hwkJlNpALcKubq0Yr77Ns7yfRCfD2xQJLVdiJ0WmnQZ7d
T9hJXN+c2g/YLfe8iRJ6O/raE7hFr1gCqXY78HPptQ9iM1ZWzOyVB48Jbie6m9SRf3S1SJL2yswh
z+JV/0tZs6gaee2eIzlfJJm0Tl/fGBmukvRLN6sKStPKMN1L9vqJfzUVMGLC7pA/INus/CZAkISV
0QaFW5+vFMWA+/0b1kRQOLnXWEQNgzt+GI/xXl4itcZmFKNenJ4sf5dBXXdkG8yKdS8gkkDkI7am
OsduU+o9YxZ+T8Zl16/MDHgBYRKdadSJ2QAqpR0P2qFad0Ol9FqDyDRt0HZqXycHdCWeyhW52DKZ
zi/qKomFPBE0sZp/qRR3PT6Z2+xJ2ncH+BNZBh7Bw7S930vfyR/F9qR9ASAqS5ceaSUF+Xwjcw4K
l3KeDrOhvyn4UuBXBjjeJjZ8t5q3H4Ux1jfhRe299DZtGmPKlt8ScKOpoC+iQM3jnICiZjlLEx9i
lB8mPdyB6l7FftTWmLl7vrDgOqSpG76G6nDUwo/PlCPpmVUsDwbJo2WHoLEL3E2lygA1J7b3+Ng9
F88+PixknLESeWlsR1aE30qwYfyxigjf8x0m9JRMYG92Q6nsdcPygDi10/NTn7Om2RpE5XzumhOZ
Bu8zfKK79l/Kk0JjHP2G5rMUl5dCSZLczzrmaFdGEaL/LjpqeXTspHRkqGrHdU58JGylyrGlUOgD
/FIl1xwvU5husP0ULK4ebvwQdOT3IF7+xvca3MyzDvsFtQG3ihj2ET0yotXxFNB39pwk3qZq1R//
Zl42Yv3KHLY5K2XSgp3Ll+WPhEzb5bbD+VHnDwP+xqd0ve2slWlxwgdL60vBKd1+k4w5KZLnQ7la
G8IKZeWHQmgarJuUMLOw733u3WN/3nX6QSb0mpgt3M8LfgC+rBtfMU6CoYnAHEV6AYz4JANiEzz9
29t4DhAX+YieNfeeBitmVnX9wVJw4P3hwSDII2W/DVNQGuOdCvUOekfVPN5Tusfw6QffSvmJXnWC
tsz8wuD1toFuHPVwYDO9NtOBK1d385EAnGSVgqliABG2ejkw6hr+3t5zKCORM4gcqoqBNbBpTSDR
5ABHXM7Tw8d0d95ign691aHDUcZbLPeXK3Sa5Y4hKfg7AsQKPGx3NyWj66BtX6Ov8n47fOlImYgV
3Sa3R1MrqJx1clEG3kkto7AoyB7q3zU08cLsa7I9+4arT5G+IySIh9odvVL5BjRMMjWmnCuTRY8c
ZLkIxhnKf+Plwju6iNPx+blx8/NvZ8/0rhAwTAT1LIHK012X9n4va6X3xQtFEbg13zNshq37/ECo
+wjnQJHpMFviHR6BRKxSA7GeCNt7hVTeVTeuTWITTRRH4IBXN487ID5zveUCE+MAe/BNFZUB4VkB
rVsp2lItbkAELquu/epEhrgqnooTqQdGSiqsf/hVOIssxkHN0cPBgV3PJqklcwObXuRGRgZ0HU1Y
fA9QiX2vdu4MEw1LnY0JhvV3OitUV6fQ8W0CiSSwGbyINzKc20RfJB9Lj4YLXVSElOlnKylqj31p
1jcAOyTtfDmTwWApxUDpdvF4km2z4q75f9sveFH0J4o4soPepkUwy3X/EwlUi1CNF1Kajh5dRtX1
1uw+OXfmpqEm7K7PhdhZs0hjuceLMG69GBguF1mnzKaaRDfA439FclTn29lb5crYZNPHDs20xstL
ijCyiWCGBdyrApSCDBrPw8ge2U9fhZK4go7JiTvKAXUjDiB2eMTE9nPVnod4XeRtIErAbGB++eXY
V2lpqvXXUT6Yiuv7pB0XCd4QRgqtex5/QQnxo5GDzcS32yvuWhyobCwRdixtoBy43ZYgZuCLZfT1
KNj9gC5RdZIiwnjFEj8NNTcRW7xAOzRhwUONqc3SxzrVx4v3XK53xJO4WWT9T45N/go3tM7Jfc3j
jrjEQNe/hVEwjUBtQ9HSqPqIpQhMoUkyovw/9MBbI97OiOe9MPrjcAW5MGchaiEO4QI6GmKLKROz
3OxNxZSwL0ReI3x76tj60cgGUeUeM24mAC/KmNtyx5CFa8kgEdDcYFbdUSsmpNTiyD/cEL0NSLfq
v10huLwv1sqVkJMjr/hw6YwndVCZRWEycz1V7vFmIhLo96VRCKmVq2IY87v02Gss++RqUXijVV2d
/ALOT0dQd6ixnk4h5bvJMflDqJPX2TxhcHPWmoAP3b+WM4z+dEDxzSwOhwfVPaJbnBgYaGF7M+44
v1Zg2qBLf3hDLg1YTDcTRD/pN1EkgVM8D6u21X4HzIhqT7LG1dhs0WWjPzdIvxkXGZjLXRVm99z6
zYy9Ymwtk9qdyHblAUAZbJMTBXh4xao8LoqV4KrR3b66SdIFxML5ro3DbpPADRAkMzD6gQFiHqSY
E7eNZlb3YfgFHuhDXQBu8V49Pr/hsllQh8As4FDBFxhn5xyJhFliSlve8k9qBSpXOhlEepe2IkKR
k9SE6oJV0RRl5okLVVyY/igVfKtPW9Q+7KkJpfM06QKPwAdZVFofF4g5Z7e91gZs5LerbGExQ78v
/gSrh16HK8WQJq6oWLM7XGZ+Qaz4WAaUzTSq02YSaJN/vpuhZRIdQaY30VcoohkBGDSDuEGV0Fqe
1ccjX1SBs/T+wjSkPMDGfPdOK40o1NeME3nR2M9vBFpkFNyLsO5Ezn+MMNm/oeNkmtZzkdxk8o1N
Pzy48AlaTRLyNUGCtj1B620/9oENlQsDb9ih90NdOLuniaXRpQfVelnnBwtU6SNwF7atVSH28K7K
re42+Qv3K2nH3ycZvGpSUW2fFQxmeWKU1VV1Ef/EKasduTjBgIBXlhzgV8RE5v2nBoQcY0LEiZS8
0VG8gMH95f+ZZFZLOYTwQYZUyFN3WVEqQAHg7zm1yvHoKaje1372V2P+lI8NesiPhuPAkovGRboK
6ByLCcEIl/vJ4YCgo8FtF2qQCIRsOAYwBxTAJzQBtHMTIzl1UTb2yGNetLl7D1NF0E0UR7mZ1ND0
NWeU17jt4uCBsEAJwlfYFWnT4Ytz5BQgND7BuTgLfjONNTE3iFt9GSmk/xA18J42RG+J6fLyYrs2
8j1WgCxtNpIe0FdOncJNz8XYZT55oE6ykZb0q3IHfc0ewmMzP+eT9DFqVb/VZYAItFYRu/oWnPAk
QQEHOjlLndNY9qRVOvzJ4+n68JOHXT+yYOyy7TluOV4NiPb+YggZhjDsUiz/yCS3Q1bWBPy7EGO0
wSCDBOqplF9cgAb/25/5KZ+Zcpdku3y5OADmRTlqLQtmVwWgVyn7InYlYYzE1DDanjxyx79pNOOy
x2kEEdfVMaX9Xstccl/u/ofRjO8Fut1yTxcpbsylXx9gDCGwhWsLA5VhyhCVB02NSwjAi5BF4/xL
SMGOMOj1myiVZBYuMl1VNTYuNx+Z/3Oa5elah0I0A3ZIpHr1np037rLYvi+m8HoboRAJfX+9dmDf
UAp3Fyc06Rjag3acN251nI4TGqaNM3SQO4fE6MoYWXwcvBwG8d/av375wqmwL8r3j+oRogCaPfnn
O7/U44zYlM6Yezjg0pBTYz+bUfkbABbpPKEcLsef6juhZfVdNIDoDbL3ttqHpJ4oBrMyTbMHcBxS
krRBZ2+d05/MkcJeFLJW3Ae0f+yZUJWnTtPEeH/Fic6F+ruACKJl70h1AH6LfAhNtrxiIuWQinjr
NZO+72cyPk0DsLyeA4skvrvj4gzeRJVmAziakP16LQ49nUnYaCcvk1IuCZV0DD2MD+GLWxpBap66
4Np94Nnsqnn1JpWdAZK3aZQTFxWR1+bSJQp2N4ASao5QZQ7DcXmIqZujzGPzQoqGSUGsBTRta4zQ
urtfcMNXwGq4cHAkrwOl857lFzsWeNU8VrSjzKywC84CH2d2rwyZi/mKBpAYRdZxQKDbTHu0x2pg
Od6K2IFJA8yjXXi+RHRjvPrytPPNxZpA0+zhlLRsXX8ALCn1yUq9pIywhHGvTBSDAlzH8CwwxhlJ
5ycmDVtmHcv7z21XOZbNjmTEcrKYPaWWT6IaozA9zTM18JuVD51YgIr+BNC38TcLk9B0vncdu6it
WUaHNPCWd5oPXZE15QzS3Svr+4E36Qf/I3cQr6ET4GqZqh3TzgpreTJ0HtNrL2JaeV3CYP9M8hRI
GK8zyNb2lEei5xLRJJox1hd9/2d+PzkSQdptOMskRl8Vb4JqfEiAV+dF+JNCrOagSaIW2XTMu+CK
JzpgN4cZIiPSLxD3ofg7Vn1+VuYdvcYsZW17Ru7j3bKGMEw1y5a7zQ38x1/wA3YAsGBwkOCsXKp0
Lxv+9o6uE2FtaVWy96xOIiMqPbAS2/ce39cTr69LGTaOVCbWo0eXPBieyUsOrvDJHvX3ElCkCcEe
OIecGrIo7JtrRdL2TSJgjZg+ObOZG6iVmeuHjufa3WMFSxCkfMxpnXkmBCh2//XGlkOKmfgzu8Xa
YHm6Stl/9+2DMm8nVCwTcIIdxSF68dEEP6SnlaTzvEaGKQZSWzD4nNrARTEjHdDxn9RXI6deIL4M
X7yaRYxLknb2yijVLXOLJ0TSvThIUZiRnkUUuEBTs0Amz5dFalYC9JdlQWdIxq7lA3sat8jHqjLO
eXFi0wJd1gGQ304xwtCNEdl1S+pU6VOFNPF5EjfEvT4M4AtYM/e2ZYxrCRcXrYEeGXqcBOzUgIyX
HJ0MD/24r2JxaUN6LJbyzWMqCCXAqKcC99V3EuALr+XfB9gMOry7nN40D+JP7A8Ux540fuw0WZWl
JlYKf0NJwC8y5d3s8qxVFd26VEGMfNpEQAA32FE4Lk3FfyAiX5NVrPlkKg6VHZ4h6e9j+2gY8zty
GzVhGhssRXQvqDTSHeWeN+lRzi5NjF2xCmVOVokl9WE5NFhRoeTQb2OnbpjQnW7Lt3HgCxHnzRmI
Smpf2FvH0tMWRxLhvThOIuzvutqzrruoW4F1wLxNudeqz9QwigaIflO4aBHol0vjoNaXFZ2o2YCL
Hze8KNl2Fb50ITYRoT9xJx//pMnUa4cJPhBi5b6Ca8u8UZkL8KIfdEipS9Wtde2A54Yee0mgYgUe
ZVZjJAeCaQ9xsd66gdWG6zrysw60GwdA6RW5q0sh/MgaVz916jqYT9+ghMrmpT31RNjp0dSCove3
3cuG9iJnE4eSoTqdTXC4SWQBcv3Wq41rPbPmeHQuro5vPjqBq0GWxcx2DWDvcVun/qBvDHCpiWaG
fRqtjMb5+GtS6k+5Lp6UOoFlrG52lI25NOqWVnfqt1odONUBy/bHJVdZIbyVRYxlH2BZusGdY5VJ
Tod71yYGBJ25jJC0kNnNsHAiXoz5ljtkTplVUSaXM8Rgajqq3AzOLU5oTBWNj+77ukmt6t/jnJBO
Ahq03OvUvuUit3SW+BtvnWC2BxyVOsZ+ueT+eA0V/TTWFFrV/LgbFwH0DMbJh2rXB0IjZyiihlo6
3z6PiFnQlxNCnXU/eEKMqprZ3yD1HCc4sgtZpqD6P3QY/NtOIrbQj1kL9D9i8cEBoOFksmz45MmA
/1IUq7ONIzby4LBXjuIUTaOj9eQYN/WjZ/N5ih11AtYOSumqSFZVQ/v1+3Lz9/xiNNlZtGEGUlZQ
dcYsls3QAvEYfU8auNORMn73rj/ikVvrUnVwHbWfFKFyUxgJYIKr1KSBQ4HZXS9S//BEIu0TqqT5
cN67y6quW+7ksPn1qKdtA9/0BBh+/1cI1JV2IP249SOk7830oCvvU3xigKtq2bi+GMuXNWQAws+8
pt0h9OsWO1Dby15eaXld/zUzLXt0V2uuZX+61OvE05x8hvJxCIEZ0s+xBmhs7+gRqgkOa3EopRdC
YDSj6RN8oMSHV5ccsaDPX5X5vOEE59t49WFJgB7+EVOLMvvpjryYYrFsPGQDpMCo0TE7UJrdLYlR
iTyWnH+KNg8fRJLE7+vi6vt7HsNXZTAlxZSRWYD/9sFdvIxxZEOM39xwm3cc2fdwsKgmiZ6t0xNF
3rA2vKL1XsBEhHszq4sTTqwYkr7XJk3SR4ca9+t0gwYDmoXlPFM/lPTvougqO8h/9bppdiNP6pRp
XCEt6KtKy4E9rGWFx9qP3jA3LjcMZ3Y+DJI/ijKs81HkBYAEFGtfgwQzEVoBcuwHKmmjv2WHdk9Y
EvA+rGGaHaZDCxrUGnvgyap7tnNg62vIgkce8eY9hRNTQ6vRTBTDgR4/AJkUYkkCBXFAyUL1enhm
98bqX2tqZ7T9p68l3UoNFkzy23T4jlwEUfuAKKSjsIoadOszwDAfSG8/eWfFU/6Z/lmSt98bABDO
1wvBd+DWJIerXIoVxe5qDMLTCnWm4gFK4lzIL/LUFRKhr0hpXCSnJ8QyFnGqFELfSZ891CT8Ocvo
C6Lapc6fg4Fm5n+jcX2oIRcmzZ42mtPxBZeNEUtqO9gnpRgM5BdzQAs0kTPTSClv43oHxDCat7pN
+G/6QNl97DCsj58AoNfQebqJg9Eam1FGq8uJ+EloU6ndH8dLdHGV9TZ8YRrfderxap7UbGpY7KCF
WPFHiutujMs/nZvBK0BdEDd83oc1WUCw+RyztooiWwZYZC+NFfJF5cPUYum7/0AHPSUv2BaWxoAi
WAkS/SEZGGguXilyCrtaGhgrq+DbwLKVRyayU55IyYMdB5BdeWLaW3E2Z30GK86Fw1KOVAyGFhYh
TEchE6jN0bAeLx0MBveYQpP80uNONBw2jutXM+WHjVt3/mEQjREkezXwxVf/Pc/oB5Y5viiBcV8f
f4cQ0iT9jYDNdIJyi15jYZSw1KAidgzzS5hxIjuCTMDrmvAoLebuMwq6pCbAXkjGwqxXLXdcHEX2
C74dRwpiWX+Ev52LoZMj7n+jHkPY5+OMcgNgSenYdG0iXIjtLU3HvDPZJeH7hHq+36eVNc7sO5PG
5MCHb1OR0RaCx0UT+NpQJYxAuL7TOW+br2m5zS+3v/JcgGz1P8ZXc8SXtTZz0EA9ukmwCzwdnvP4
MHeL+IZ/XSD8yDDNj/cdOusBJrj2sAmRPlojBUbddpv/yfQq1+SuX4uUuB/YdV9AfTCiJURffF3n
2KIPQKW/bdqCx8po3eWQJSNaUgjB42ZMME4zFMErK2IIPLltAULfZMH/gFIzAsdYd5uCXBJEaHPo
5pRmqJb/uPcY4nFac3XmWLTXrAho4Tep26M92H1GdlhEKi271mIJf4BgC+VsxGhdVqJsLTIm9qWl
lTzkYyV75wrBktXyvwzo8NB9393A0ALcsDJxWEivXBy7VshCCioUw2STQVsPgdO7l02q1nqrY1Zq
3CvO/IoKoJBDunVQan1GXNgp1VxC++JHpSfT1plZKX34CSgQXsvdWlDzMo5ads9ez+BaI/VW4HOw
EdDJFTVBXExc5NaxTSb0eUKNObUHC/JdVbHxQQIKw9Qa2/eka+Ic5oDdFe0NFkVDXPF4x0HccOi2
RqjbmoEgxNBlYxqchTDwrHcNhFl9pjyEG6BWOFBrCN6NFQeDyQlSwba8/HEFIimzC6n5Gw8UqUS8
DUoIyOyUTsqUSeG0TLcYkx/5xOrLrg/tVkkSWDiwo0OVlWBDIRnKB19jzWV5NUfTUMlS/+l0/Ab4
ZsMMenfLNeU+Drj9ozt4t+f81QENmkXoyVEW523DDyef5+CWhaMVDnHUFlM/PuzdtraGRnoOEgNE
1k65YJg6eCghCTFhxrhk8HoTwO887FJvfpoBpnQWFa7sfsud25j2VoXBNVWbp3GZ4fA8fsiy3rLv
AJi+bgAHqNRYeGg3l/hPKlDd+rwUqAfXuVwt+JRvISQdsyDpgN8vsLjlccUDuXuZF5mBjwEnYhg/
UimRUOiKz8ogYsgVp7SQI2LhuO6tKcApqgr/bNkWLdoXXGSl3BBiUZbVO8pjHcF9hFpq+DAYl4Uc
9K20k+QNYFngQigMlJGGaMcEdp5kHg+340hDRBUDu14D3n7mHIZdqhxGS1BR34AV0HG9PB1zihaF
QdFIGcqX5WOYHXfTsg0fnfPSf5BX2jrkHxpyIWeqrXSYZJcFjSQS0PtHm1GaUbrzToKXsppsIE88
LbVhVJHqiemCAv+Z/opcZz63ZkBRmVltamIkGLMqzBk5WWearhw8adfW00eraH/KJKwwl4ZkWbKn
2jshCvQd5qb4u7lCydwRv790bYEkRmB6AZHNP5kB1BS+kb4/hSUJMu1iwp0UCrrSFyky++sF0k73
2Ot/KCq87YRemY8TTp10asTKOTULGChZsiVNprr0/8lQoGlPzUWe3dgIXt439zZcM2zVrK94n4Hm
mmiYGpE0Q3Bv7bmhJ10WYHFpviaqSsIcYsHXlaODIRaa0H+ib4S0Lxbp+ZaOh/IgjA4vwbdoBYCF
Lqx+pdOV+3mQTDyt7jsSr5oArxxSOFpBeQSilWtGxmaqXQOJirLNWhbGey7XKNwtRraSGkl+OLsP
5DM0UqE3oKSKurJ4yCVCtlX72VAobTLOWtUfdTab9QOr55KLxiLE6xsM9mGa7daJ5bULU6hLewEX
CRk5zCVH6jGN0H+0dUCG0ebs1CRIzaejyzKBEiMwUupsUTtsOOIS50bqho1WGvIIHVIKbGN4WebR
KcbCx3O5l2tmxcLp7Hd6q29vnxxKguiFi/bGUxQmkk6vlKlP8wXNETKC6SmB5QYiAA0jEZjaUOzd
G8uMdmaMyvCqp11LZB0uEJP068ylSykds29EoT93/yEV7KvU3WVX+HPp1lIk4sCpPSPg4HJkWh07
smp085dCCQiSXIOCpla9UW+Jr4N1IlVfgba/62JMYpB0nx2fx0q1IA8Tnf+z0t4DlMOGUr4UhIvy
cDc3CLyyui5Oyt1OR+d7tbMWNVOdKzILHOISwsQTUdHIPRkWaNp4SKZXnKyOZwsp9r1yIsJBv6+O
Hqc8F1zGRwx9mRARoFUMQMw7dvAOJ92Ytbb5E6yhIsP9cYns3pH94RJ5AfH9Aaq/0wqKQoySjjM9
ZyIq16iK7+fQmPPuMFbmmAkSXciNcPAuVUxTvdokl5DmWP+YFl2RCKJOVKzebt6iaQRo1y8vipRU
iQs8ft+03oqZLynF0bXn0eSUc933D4u00Yz6gqIW3PDkbXeIcl6w+8SzhnWWOZX6XYjrl3RCvacW
rqbw7YRfUt5BaxtzJxfBUZGJ575shMReFoiVKId2V6zfJYPQ1+qUrIyOXgZzNDmH+gHbjrYX68za
xC1SIvcUXE3DXRyYiqycpwbW2PaoUOXIRLh8+pRhFiVBRnKUDGv9Oy8zGOdfSREXOP5va38DNg2F
pZs8VBMmzdqBcfxFMJHnk5LR+aK3WKbDHW9D8cMlKJf/3P1a+2/7ceys7gGYCfsTGNZGzFC7dsaj
J6ZpEID8CsOnCTV/pBqbdVqr0ZpW+PviuTtkEpPQpoJdIcFhL3ycz9sso7CXZBpcWwqHL8t7jdpM
Lxx9yymm9Hc1jvmb7qOkNDOFIWX06347Yhaax2wC67Oky16oZoGwACN2citjn5QWxWkeAGJgPp/r
3uJ9j2j/bTfNX7Tsmv8TycNGJCq7FDXeAOgTSPHW0pr+wlhq7/hdp9Q4/d4z2YHLoWXn4ZZTZBK+
VVL+eOoQgZOE+y1xtSsKWlNUVLWCQXAz/x/dBbw8h7TJmpfLL2uphIUSgna7jgYQAuHNV4KEUwaw
HDlh7pGhSEGlgm1zBZGgxbUb87kdy2Jx5FVIihECXo2rsC+EYUInHAJSAD1+rdqJm4BIFLziy9pe
zZmy2VaVOa6tD2hq6raq7sVWLcf2upbkIusVl/AlsqjyrHAy6rXOgK29PqCiToZoW+T3IfT//Sij
aPfZVenJ5FyG75TVOBFb5n0HvrYSsCEcSxM42w3K1hRzQpsK37wBkOnoqiEUtBvE1ibKz9H/dr7+
bONsyJcYP8wXz4WYbvaYO0sJjimX7oReiQKE50c+5itRAdaUOgPEz2+7kA5MgeUa8c+dzSkypdR/
nCrlTt8mXOpiWNhNfv6QPIET+3ipM6z/KH3EatbVaBIwA2WviJO/94lTGF+AA0XMNWMJAms2Mj3E
1jSBtxsBPna5ig2KCNUszXR1gEWdy0AwEQzzf2cBKcjNIbNS8zlAD289q+ZY71FORTFPRevUVhjb
CbJp28HRW+9vMhU8DJN1CWxCiEjAnBciCvKqrxHICLQvI4Mk1VzzmJZ//dUKLt3RhbTGjJCxKWWV
HQTXl+5MGTj5EY0ApSbK/R5I69YpBEvIx1VlnD/IOXDfY+tIts77rmODe/k/ASO8uaVkZUuGW3il
EPHsDXdynWLNT3M18PljST56aMCNrte1giWnq0lh/j35T0PV4a3SJ8QrJcrlZ097zZ611M6g+3PY
mrg1k7LOo2gv63Two4uUNqEfCAr2JWcXHNDaMijYZ2374P4CDFXvo26Ervi3GTxmjjhYimxHfc4c
LIXweyXn+1FtdTjSDMhA6KjReZvVFi9m9RPncc6khS+LJh8xIdtPFv0muNJEouZXyzFL23H2awOh
f2LLLJaJ/r3UMr38VUkQkCyT8btfy+SLoTcYzmA3sBx1eu7THHtkKJvntWhdBAjRbwP2ZOX0KMyI
V3LDnXUxuTUz7MTHIeVEJwv5hvdbsvKMlWBmI51wxNt1KZXF9ZLap8wSIBfEsh9z1Sfelm4uMEw9
RVRnQqKc/4oFCVfVmU5H24M2arD89z62r0Q3CNTO3xqVNMSIuID95m6UUHVWG/tyohueCqJnCdf0
cNo0Hrq4VgxcYmLojM6smkEsi9QaygTElYjX6a7TGpjzzF9nV8n+fltMJO6NVGuBN82mBby7P1Gb
ByS9MCw5nkQLhpwMG+eW4JSsH20YgRNWNXO/H5tV0JFXe+EotpknQJNbhdeEcqYe9LB/weCeBu8O
hnoJgUQy9pITVemvxlLAM2o3tXipPhW47bGCJz3KahxiLqbvMNvh4/3O0DxA6Hb5Bnn1dfu+LxJ8
HbazSCMRUovHYuSekClpv5ObGmP+885vU/L6P0gpEJS80VuyO7r0OYh50+Mkm5kNchoOOT3UjiJw
8DzUleCidEgSlQFcUDEb8oJaD3OW/x8i79oN4hQL2ftwzf8BQBI/CKRrtnMkjl5Nzd1UIq+b5Tzb
anix92tNQ9r3D/E/mJoVIyXYRh0zuSfVVSOPB/5JrRn8h9R51cFAd73pJPCUo0NqDtwfjmhbV+ba
QRKLd4aSFJOB+IK8HUGXJOou8za9t8FXeRoM8dSybWf9Y296L/gGoQt9gK7zKBhNb7qB6tHLk6QG
272Q1EVQsWS7jcDb+zmGdpnkHZd4FjEUmBQYNjPAw6i1h0gF+JEuNq39xwCnEp03wQmMx+FWJfGf
Nkk+Gx5py4gwJSQG2742tzF0Uj+V9S8xHSL5iHAFZd//q9rH6p6bWFM1I0XC8W2F7gKD/wPk4QlT
CbvgmasfkvS3YyA/pk6v+u0bZFosLS5BVNdHgq/evBFjvk1N9wjZzRkJx+8tX2bOwiJLygjs14S+
TGfAGrAQykd7lI8j964aNyzqkRC8bC3o8TpERqYIbAHMFBLXn8OeNzgd/hwd73Is+GRGzzZ+9wId
XpBEWWqf3j/jsd/+Laqm/aNWArKid8jfzrR+F3tLApU2S3L+vQFNrU121ps0V/AyWrN5mjp0rFlp
XrDVcUJw25gzwieMQC5Jr0mxZrKTo5GP6lmtmLq79k8U9v+OIpEy340aLJHMQBY+Psf1t2JllCfG
ftGEvL91+VRHvSZ63uJASneiE3Oyu2fB9exkAwSb0qEY7waRrMDo/VaRQM8OJPy9xdVB7ET7ft1v
zHuSYSjn/ApF0lbRbD0/WMVUMI13PqKGdPi1sLf/axn0ER9EBnHJ6m3mzoDaHoI4h+XwCs9726fv
2Zslc765JNIApnKdKZNWNkyHCHFLTQ1wfO4fZd9S0XHDpxfa1A1VE2VrOUNWsCYuboGcuzzCgR9V
JRxYZ1TLsdWq6O8U/n3Y7z59u4+GeSasBTB0f+E3u0yVMJHYMHzbWeKzCere5SoQhXWzR+7JRluN
KDEADc+5pVv8/3RkTVoVl2tnOg3kVT2yt0icyUwUziMEc4NfWJ5Rtanwti0iv0ghing9f3Zq4cpq
M24Pm+wz8ktr7hauwmV+dND2dAo2YuuO2xqJ+bePFzUDKCmzR5ikKOsbDxVpP4wCog5iZM0k0hBF
CKhKL0zBbtZlViKscBBzBZCRSGqILdnHUpHJCqU7z5SdoKVp65F8cNQBwrHnhPFK06V2qdAAujr5
00wufVBhKZv09v81zoI0PUSGe37XpyiitXvrd0EwdQutFCQquaqyJ+756JQt9ltAEF4lUYdHGRXp
sUa81RtW84v7iPzKEHkXKabkaQ8YuFUgMUJNxbDn+WCaQPJXwbxF+YK+qiBzyigjRoGJ5M0PDOAr
2BXST/ItanRMGLz1sC39lWcX6btIFRKZi7Icg4DdBYyLrvLsfJwWSshmXxOtn44QqD4eZMgvvuwB
fHNmONRA8iXwY3u+ERy9EbsC7CMVHM3n1Oi4s8gvwh1XDsz4hLF6B75BE+FYGHaGlnNBZY7+5ea6
S8kb8N7TyP7lxI2K3y9Tw8q1uyJStWLgyhN4l+XhPjgxKw1i9sxcXfNsh8BcxFdtCr7uQlf4Q8mS
wPMRP7ngPPL47Rl7fPv7RGHpYsGHHYZ7PVBUoJBm+uCEUbJbngb5kRJCJCwazAQByt6RMep4w38a
h1F0FgA4QlA3wYuzoFTEXSA1YAZF5sjziSK6/yDJGphFUN8fCo8AsWBvLkcZv6400g3/0N8K88km
uHESf1E6LB8yXXCmo5xjhs5aYvnlODPMPKTn2RcjlqgTKuuoIOGP+oDTwBh6VRMG7ffpV9mNoDN0
d5hnX5xJMY3OUhHQ7P4nwfZy90EYs75NcNyQXO45NnI1WsqxVSgxxdJIvtA+53fgMfHe0vr0iRJB
dg+AzfpN2Om3nun5eqRV30MwxRJ3NfteOPSBFSM6yCQed2/ohT0NzZy+eTwpDMwhqHM+APJiPnLG
uLET99Il8gbAVb4/P7DOeP74B4SSMUiD/se8yvxZNVmWSDvSdZYVepvzTd2L0FwqCi18Z6oiRblq
qY/bw1q6xQgwVz11PoetbtdfDvXRs4ClUhx1YJ4tgl7ilAMq9wuDanqGjciCj06VkM1AyujumhAT
mqUcN7b5BJi/HgkcL0obwBSBJGAQR8IiXYH+HCXiSxwwGf3hkUgIjRO/+XamqqCOCWaqsK6j7PMT
3wKVPbzBsS4L/8lmxmEdYQJ5McJ8sXtIY6Yup0K3UU2rFCt+0UWZmJRt1AVAdEHOzWcCYYGg8b4+
CmCc+l6rwOdMjdy9oDcq1ZSKGcBitZHbThIR+0rwmDN5kK7DNuovOSg8GB7VEpiF8yD8XzCyu2Pk
ZyLqQWSB9NxgSycfpBceaWLpvmD+s9JTU16vPetYDFGN33tYblFWsrl/VLdZ0dCOhvG1pbdG2qVT
9aGd8yOw/yfeRNIrF/rMneZJbDziIbZ/NaPCLAGHui4yRFxd3f0fZqLn+JveKxjazVleEbv/jh3E
YKLh0kkVIvuJhcCGioUDFj2Kllq5qFd2H6cDBjtFWjjZbAW1Wycl1wFarS35sq80ZbnGXp90r0Cz
Eh7fOqntNpn6uHokC2c1nS3XSKgsoEi6OwoYZgVmzA6M717VRHT3iEV+cSkS3aBuaNsJAIkeFC7n
zJIAQwMF9QLQZlExRvxmkTgArp+tQvfudqD0g07SqmhiFpFPt/ystoei6SEmpzfzP9ognEBdMvFK
/wMz2oYHPBuBra402UwOqIdI/Y0FOXX3mY9Npn0hlYbfPCmsRhBSsY3RyG0EeuPP0F+Mh8Cw2Cf/
qkwa0DwfZNCGy/XmdxQ2bU7D/JQxz2/0kZ54G2aPiylKTr7k1+BLnKBB61kdM8x3AnoUEOEh1E5Y
IjQ2uDY6+Ln8OaAxWQnl5CZvu5SBDDkpLgRkjoXhccGkfQGykrbvnTtvgtBHZ3cm1tJYd5v8xvVh
py++7IVxOkbnHfH9ml68pJ7b7S+/doN+OckMoBA47yNw8O9MW+dgmhMUdC/P9Wr9K8ZCFvpydBcD
lbJMBA/J9RfVFb7U73VkJhIcd24nEF4is2AlhojIT405UR58U3iyu/eUAVwK//+Nm/nNxuuuFNGS
fExgtZneHO09f6g6vflVRhDze6N3dWULIgb8g65DH/jPS5gyvpZ2T0ddlIO1rB+guwJ2s9EUa7QQ
zstmVPq+BxtHDfqJc6N6BIEClQfzDkpSlMyGPHNhIpm2gk0/vXXXFhF2quWFUau8RiHfHYUxP5I0
lhXRWY0RTnFQsJoOql4B+z+c3EtLpcaRco4AoW79+40Ya+d0KkuglcTvSSKK9iGmeXykUgypA6XZ
DLVP6oKhzbsKB+1g2mJm1WJHuwkhFzHDDMTQwY3Fb8kKIvWHv+nSbwFwOJwDw9sVTR2qdp4w6SbG
H21kGQERDLoFygZwT0i9r6gzY3Sy7oljVaWEhBrpvH8PBh1QM5LCNCSfTAAvuW7Uk7rt5kczh3Iw
fTDRnwpGpFIzBn4v78dHE6pjJgVbjI2UUno4FXirhdylVTmZnpRdVfZr6Xf6FEXyxR6XDO5SLQS6
8+pz/YIQOEIbKkP6RNM9K7YhLD2gTku327lp3ZJBc2V6o0jvP39PIDA0i83347Ihf3ApY3TQzxsp
naxS2lJmWuL80RxLDl/R5QUixBvrf5gmrEXW/qgY8rt1XZNjIk5OqmgJhQtJzQ8KqiibKHkl0N0m
8LsN2YbY8d2j9scu6gn3e88UwNfcA4FDPUQ9GUnpEbewj0Pl9YcpzsLuZ4BLOU+qPGFUWTynpJtU
d4zA1ziyolcb70DtLH7mn/Dg/gwOTbX8tPE0S6EGltDPe7DKu/W0lSR0+uXFWEcQFB5PTNpZHJQ/
2UkzSyysw7KrQB+gj5wwkC+rQgKAmiMCA5Jpd6kBZ8xR+YsoDKC0fs7w3ahWwcz1h1X+iqqQy1Xz
Dh+FABeuPAwB57L5YnYtxLXOLmZJzdHmeZpXt2vqyN+YUo5dFWU68lgnCxlaAlI/Lhd/qSUV/Uzv
BvvAIgKVMLtN3eEpctupWestL43sNX6d5LAmePUA3o/WOQAS90OCweTCa6LYSHqEcnNa6n4D8e5l
4n47WGl5tBIXKmkZMdJ0fWde5GFakVVyTHjJaMUxSiYnBQNAa7EnJNjtyYTDNSu3gUxlGC1jrsWJ
oQsZgzVddRVqRpgvGHEcrIt1r7t2vfUQyiCPBXBD7BZrh91zUvhnnut4puLbk9Fui+z/dKU/zPDH
n4ZJK0QiwgdFO7xf0cP6Uf5cpd9E/LPe2rfVzddFT9wUg0ZstizpBpeRcI5dU+wUtuZGEtIL4g1/
oHC/XrCrDNvSPSYolYHYpY9ykOd/563nBZDmTwSNBs+dQkb1a3eqzx02YxlEOzJ7HCqf8Eaqfn1a
KnggPO7ZxoHYq1kx1z+ke7jLj0JhS2dNOJ/Ddr8xaM2Zv+Gn7dQabMaCEzzcgHmxMHhIxe8mIkJ5
IUfuJuXdJOxozroTtHC3TJC9SmWMoRKF5xZeEkrkKsO6jC06yuXkDItF1Q2EKXyX2tG76rG8Nd7s
5bzY3oyoswBkKkh71dFruTktM7Hzv50pGnm0XVaUXUB/DdVjL8vJL1STijz0oc1mB3ekeYqheFLI
H/oBsuATWY3ST0RmoH7dgVSExufX9kcOQ33qKM3ba5SuE6qE3F/BpQjHvE0DJpyQxSkRvdgFd/a8
dsr5c/zEstFbe/mCfeIVITtZO4qp+uK/ffOB/0F6zp/ldFmCAHrBNYyi/BgWh39GXEazeMqhtkfp
6R8o06Y8w7OAuosnti4x9Stn1UNTXYZtHwKWal1PGgyzQmAazMZqpGx9f3QwYr4cJgjRlVP8VcdK
Hb1HFE7+VeI44r1YdgCJHnkO+LtO0jjlFurJbvA3ljbt5dm9AGrm/2uCpcFswbF2xlXxKoYxBL4B
jMuCjEDDWKZk6hTBwZwT9bYWMGPAC2tRIksuDr9lou+0ea28Eq7C/B9PmCgHfDCA6KmfluoALXE5
MUJbGLDr4KOnzRuOPjLqGi3tWKIqf9h0O6Dk7Xx3ENKP/NtI035cVmnYXrXvkZHXtWIEtIjGDza/
ERmEXFZ6/nRazO2VuzvPNqflDheoSf7AxZLHF6AwffsoX5yKKNvAOQHTbd3pCdwVjuExMGNyM8IT
srHl0sE00DY3kUU86+6T4rhfiYslXhon2Iv5XQAx3AUUTyME/VKg3fLw6XmE1WqnslMkPqdhELCM
cN6bBR7QIC48sUdsrPC2WA+BFb3qEaig3j4uX0RmVySloFGNSXL6ZLZplO1hzHmv96wvmzSO9b+8
aUJ8YdZ5KTCl0cC4c2ohzOP2q8ClKpZXXAqwlFnp+vmqhs0XjBV4bNknH1hEO8JJjChbaWG1Vy/x
yvg/C3Cb3Gll7jCg66P0DVNpZGM30sB6kkxP/S4NtiGcH6JIY5ArYu0llU4mQVHrfddI9Yb/4J98
E5WOfIAQ8XkhtXpww5B+i9+iL2BwaUlCo3L0/p7kUN1iM8sBjm4Oi1fu/Q31+s5eD2K1va6tM0Rq
2YlDQmpID8KHlXaIpyZXi9nJ2UsStRCR4dKEmsSWGO5IxYb6HY6m3he0e9deqImnBj1PO5wuPwUi
qGYbxSC2eJdV4VQ3ttwLiphoi4O+7DdQ1RcLG4dUNHbFFuMDo2CEW/EmTCd+5QBQ7m46p7XRzI3l
4Xs90GmidGFjTG6Ur/gl4N7aPsI5H0/FCxqjeUSIniQN0JU4OxOyyVAQEsLJos7A74gCefo8FazT
yF0f4KuY7pi8SVlFCAviL2sIODnQTLzIkZA8n91eELBJEY7XODS4rdacanDt7LmPweY5VG3148xb
w0L+2X2gon+5LWMJ5ZC2wSWishdeeAN/QXKaXO3arUwBvdsEfv/QzPMmH7W786H/BziUD089yGnD
Y2P4b6wFGWiczQXZy2PAH+WQvx2aA2mVApk9cZBluwQ8MBrWmh8V67sBF+Ji9oHhuo9FPN+lGcSq
w8lOjeTyFeLI+db7EFg747yVzZ5V4cYTkOrzKDKLjXTs2XJZS9QQxgeVkYI/DHKhx21gtTbJPyJO
A1efqrLU8e3ySB+O/+K1WpCuj+6rVp4DN9zNjxVVO3puv8ezji3OZ0Za87UtJXGKbjVyRNgParTy
Y+eDBzClgbFCoQLgM4XEhOstKKEanzFo/SDBS7rj5rV+bAgBTWM0/yH++UrmlZcptFAOi8y9Eswk
KNb1iQv+PSXxVm9dWrwwUVsE0NMrwDCrzzMiB35Pj4CNV01A7eT3HExSy+dRkI2XYKHLnrTR1mGg
30aXyJ3U0DG8rHNlCNLQ69BH1BKipDyKN9vRxO5E3wpNomAgygGnugERLHyMYqv+ek1Esdj11rxC
kRIBXKxearW72jSQ3sQvbLaR08WtoxCqN5cd18N8p0ydC4tP+huQO0sGn5/grNVgIFf+T2iBG3l5
8QECQ00swiMaYrwGFExZXqeIAFveRFJJ+aSL3y5DhnsSmNdj4seL+6uEikzbUbEffvY4bbaeu5Sr
CtcgqRmuTP9lR3tC+DnQCNbWebxSHzYky3E/6KxD39R6+HL9B/vTmd2o9RFWWXYX6QICiiWkKlJw
471ct3aB9974oz2zDll6Dq1ZHbohS4LDP4mx0S0xIOJCCusptvTjb1g3lwADa5YUc1+YXtZvVc/F
J33RoLAT6lWb9FIqF3vF2Wn5zalAXnCr6yxHyaf7xaVd6oRNoYXOcyfRAw26i0LtNbFu2aXsE4If
0qObewguD++7zh9H+DhP1EhT73kTO8krczpTKyPTEdrrarEQ7EyyWzMftisw+ezkSaqV1JAgXNQI
bA6zz4FVNJ03uW0LPDahd77CLFrTrVQDqS9wiABd5xadKtm+jd4bjBm3ziI/2J630EeGihiUvehS
cag6UusBO+k3fLUg2fBKKppZvS+2chMtXDdbjhree8mFZlPtkfgXKctW3V160r1NGjR5G1dutuLk
TWQoPftopMJh1h+N4ZQWiB61XQncQnZRMTyjCu5XQNNjsJJJuuvwcP0ApMmE6Gtb2iEHniieu4VM
i6w9OWIsPdju8F48xIRywAnJW9EApZJm45ANQCDHH+0PhMjcxLfxP53HtMBfvzmPvNj96lx+1DRD
sVPMpbMP1Y6iaA/d1wP4K9Glvp59OWdz7L5qClh1h1ly9gWE86v1L5oNens7zEnN1LZSvdqsNNOF
ttHvPJYnuWEgZlOCqD3aAcKGQGPh/rcm+6vGGcAlu5jZDhg+H+1ElO3XwK9czEOvl3Iitl++bxlb
QH7x/furykhJAlrBJFJNvcGWwwLsMgVLV8GB9bgXH8sGIiTxb6cbxPLwh2FsK2fxAG6ElM1/DB31
GMeZl0IwyMMSnzzZ3xeg9eH5pSmAmu5RHF5uUmZQO2KGO4OOACQ6IoPir8bnGPMI3SuE7EJ3qltj
6b2oRWFWRuKAUca2yUbai2rhyRJxHp4DmPmmXqA+L2lR2P68EsyR8mkGj6UXV5EaYA7Dizr9pEfq
gq6iQmxl4RR8sgjDR3mKzqq+9YWq4pxZDRhLm9WxAVZWvsCu6mIm2BHbaqCVKXfVicdytllAPdTW
ZhxP7x+74BPfN4u4XBzC9Ds0EB6SM8xoV0tCe3KqFKfb5jq0F5noKUZ4e+1qIEeZXPfm4x56mpIO
dwxpHeAZXc6Gs3nWRGF870Kz1UUQ0eMydFBH3D0/P3A2UxOzOrvOIZ+t1VjrLfKdV8ubPJ+fEIii
v8/r6ZdoRHbslOf966yyPsGGiCFqJsAcnt880xjgHUv+fuvqEh7cMnSjX6/CBmxdw6de/jn1AFpe
ZwMMdRk7ksIy1XIi5eJmQbQwfzX0oWDJ12PuV+1XnraZDQ0vpuSZvrS+Mk0SCySiSbsy3ARiwFiB
5p6wrW8fwVaDTPPAuN61CNzsSsnbFJLqaeyvcZq0Sptu/R7bQhJgT0mylQkbKXwagMa7VbDWGLN0
5I/b5L74pl4X94FMcpxNMxyRzgEonpGibPLsD0t78PXQwfwRfQQ/mE+5jCJpCPHuMNCa40zrrO53
sMI3TORWtRme5QWMrtBSIz2Jn2L2ZB4pRhyzKXvjy2t5DovzDk/aApnlrTEkKFo6q+WjweZbj2E4
TXwDoq8TdIKpo6t+VDCbPAcKp2UoJAXTUmTRx43kiCqK/KLlcj/rPiDz/RMjkon5In139grhrTcd
Kz1pjp1q6UvJmrWuMm2NX+HjqueYWy8XlAvb6HeRVclAGkW/Oo9UJbKJ30mRYA3vbqI4qAi9sPLD
QVbMeUOnZQj9CO3R4pAMPnusvC2FCdj3cnyfhhA+V3YOp7KxrlHQR1g+V3KQ0RLwHGfhNTXp7HNW
tx8Qxgs+EZNq+9DqVLQmn5+UhC53b+vNOMWTL6QU+PMEgVodIb0OFH16idq/nnaOcOxJMEdXNQ35
kHfEN+U603C43RpboVaLErZEgRYRDGq8dmTPU8orm+tqWExtfxvTSuRQo4KGupEv2gxmzy8/EW7s
paAlK48ZyYxLCU7xJlX98DXoXo2ec6SbNvj/OS4lQKCD9NsXozh3sy+nB6q/abURiapUQEtCqaS7
yyaQRNbtsLITHCsEXSwMofhbHPxwGsxFnE4D/9cWTU3VwXMuZemsBGOxfKKhrxlpMWGcAX+iDAvO
V2h+ImsQTCkt7A/i6r0fSnGsvW93bz2zfHLNewOCRx5a6Y/ctsgb3ddQ2ymEHTQvdJudfAW6otmN
SSMaKWSHVZz2emPwVsKDoysMZ+tDCe1qQb2cWWiDBWZtekzAZxNMYk9VsoqOxn3vk6mfDbvjPT8H
iH7VvPq7vlIAuh6C9sVZj/X9PzurffK7CPkuZekKvjB9gjgINQd6+BuzxdZaT6eTYML7EWdhQMpk
xGknwq8SOY/Dqpy/U6/CP+LOfhkufB5b5FyXEu/qEHlku/nl1HVoZyNXm5W939ct1ARBDT9skUB3
HdYadgwq29Qt3xVMLIGvFGkvR/OwZepGvAqdQkCabRfYql2njD9K1Byd2lljFau2JnZnJOUib+Tb
6yt12pXIEDCvIvr4E5qo5vLWtkJ7VZoFNQVpW2TfEP9IEKthaNRRolgndo5ocksyD34l69NWFt9Y
xuYQ0JCZWTEjKf8k8g2stmH8J16dNkh7gdxcAl5uUArB+xaAhJ2JuVaf2dPGUZufOhOtNfdda3eJ
VMhi+CKTXQb0bGtn/olu2hwe2pa2wKjtTITPxN0SAIQRuWxhDlY1cwxVfh0fKxzL2UXyflxf13PK
UwKhKlxNuuTEfP9ZdJc5vAyO8XpUF1BPIvuJ9NghaIgrgodkYR9hRTkYc/8YkDbBXNh9O0CAnGWz
O3oOuin67nYwFhkeE7cE75G7tH5Cj1dV4amUAba38ZyzbXzx7UI6NR0F0m37/qhhMK+ru+GyFt21
KL+zm4gRiP3yjHzG9gnx0tx+HEeoV8FxhHxfMmjdxFIbceKt4o2kwju73wEh+RbJIohcao1boAr8
EgIIeJFjGdh/mbb/6ZVn7f4lD+9gPi4RSiVCP/SrXWxwes1gqLa3m+uzvpayrSzrLFdN+5VI7Sw3
SZvVbbg5HLh0oioipytaQ3w6phX7UlWYkInRrr21PRQsOBqtq9FbP3kbfCza2c/916F0UoOQmmtW
OlEPTtGu8q9DpzcDMzso1wDxGpJylu863iSZIDaK4Mi2eGm2CrK4HXrcN19s4ROY3vltoYhatIbn
civwF8cTkCmnltN6X8PwOcF6p/rfR8SORSRIO5cYB6CBrXCXWtXsiOZTP07Esg8TvvKehtNUgMzX
Bmz8Nhas10izyFiBpiK7tN/glGN7UYM9vAvQVwhl5qy6ExA2Q1iZH+7mwv7UHpKJ/uu8/d4o2O5f
5dnuWFMnBpKX001uWC3qE1DMjF4/nGSPsCdfXZiqvBX8+16cd3Z8IWAKHqNSED9CuKU/eHx4j5Xw
iBKUMsjjfKkP+JTcrRTs3L5AgM1YA05FYG2cx0kJw0y5Yh9uxy3RuYVxq9C6HN7sxpMI6F3ZiwcC
wIkLhPC5YQ292uVWNuHExooCtBdu0zWkLD/JSXHBLxcnbXFxKHW7jTyShej0xuTnKHn82JZbluwb
HiisXO+MSGQ+mw5ySeMRJF8VZhXXMv7jNR9yBB7u5KI26J7WbatSQKjmhX52+/XwsnS5ugx/Hq+f
UJWU2ZNNhdDzeunDTils53uQnyQjuRTXUQuoOLJjnph0c95CqYaiEnQ8SlxNBS6+PO7JXHqvh7Tp
W5hzpRaR67fZ1xFjh/8in6McjqN8/lZ+sQi3GUIJxE12gAvjNjDfQBW+81Ga96WyLsdwS06Wm4YD
ot5/UThtb7X+WXUDOuu6LeFM7PotPxnH7R1v9esYK+kjOs49rhxhHljsE71/jWL0yYUy2z72O0dy
cd0cChFTKdnffLn82P4v3QqqI0q28B9lYqs6fb+feN7QCH5IktLm0jy4fqS7ugS0bQWsgF5GzvQp
K9ZOPC3e5ofzUWcwP+qenZ/mtKH3o5AJkBtu8rqCuu2wK/My2WpbFAX8m0+x9zhlET9LrovGHoAw
R1OgdSOVAsZfzOk3fYMaoE3BWL8z/mla24x6YAyXharSFK4csQbfXBtdn3ERVy1Ixra1MgkjQIrf
DQMQBm/InRVA2LggQbGkyahYNhffa9fU+Uu6RY+/+h5YR+CFwd846zdillcWpdBuH4MriboD7teQ
HYjN8TC0JPMf1I0rrlvqRmfoGT87JXTk/VPusxh9CfmpN51XY+T1oQEEr20ZnUNORpE05JYTYfB0
mlxXNhY4FMXvgvhv9YQgRgSjpJuF36r/vPiQyNFLp8Iag0IdRhjgPndDtIvWqXD9zDSdl6o9nv73
AJ+EB7hjCqp0B0Mm9OYIe25K8yPxPTfk4theJB5pTU8uTiLsdAL6OMGlt8eGRtv+ykix4HlrHKNO
PhQcEXWID+YQ49eR8G2fR/of1hwdjuQm6YygGKrBLs50gdCT4aGPpCxM2nN1PPVAdKoZA0YeiQq0
eDVPe78yCY1RvE7uS3zmEx5TKdVG/i180dPWIadQ7lkBz+Jnwgv8Ch7spJtCWa1oCOYww8yR8saS
PQrAWutMcKNXfDl8KEAqDpvju9ZYgFMhT9tdtyl39kyohFjOB0OWv+q2zONjvTDXtf0cQLwDDtIV
e1MM3fA/OuN76zChgCkGtxwFWFlWqbGkHwXFdk9TsH1i1wZ7pHS5Ezr9kYngf3qF8+jG7h4FKLKU
3ZKZH42r2GiGfEpt8WFOxrjjdEJ9XhCF0E+BoH+Q6GtYo03CvrlLCi89hkCf6A/m3yfVw9jJ1/MN
Li0mGwcSBlbgLNZBeBX5mfv9s1F2XxffRppYCv+kDxn/vmM6ccMzO/3bSwBg11kQfemE5eGCuiFP
32gnW8SM1nIZG/P3CYmIcIm0vP92/5cZa7cduoMbsLUlxqjNHMx0OAD+/UbkU/1kIaV9fHyoaic3
RPMClYXUQVrKDY/OqZH6IgrLzDaTTRIrqlKrGmGPpO7L/i1b4n+ieFjb2RQJJbMfVGlQgZyMN8bX
bWDjZy9Ic0s7eYiGKkR8i8JywOSkw4L5lgdrlOoTxHUYiS2BB8W5uo1Uir+rTwnrM8tym5+Dg9Ib
7LiqX3ne91hw9zwHOW7zmfBkQSjANDeVSU3V9X3zd6ga7tCmSoR0gdSap48ClT8Y62bdJLo605sv
NLCXHypro3PbPkGZ/bQO9ze84WwKczsRzPbVs9a6jv5KOb+AhGLnaGD8vdxZWMBt+iBC2diLxNHt
ZJF0/27VQhwMkx0ED6z9eQOYbrC4V3ovYPhOycEUDo1yHTRoKQuLh0RilCmFar8+Ij9uAxdc6FMI
FNiPTP0WfkNf80+hohqPk2q+geSRTPa874VKxtZ/fXDFIg+PSxMAxT9p78vZ1353yC20zM2p/Cv0
upw8XhconeTprDGqm49j8+0OP2umyRMfhTtp+hPdkwcKQZPonVlb5VhPh79lEy0n8gPOkK8b7wBa
75nlCqJzuRDddr0IgjaFKAgPO25itqOzdxiZuZQ5EMsAJgP/1GMNJ5F06CaH5ZA+DWP93jh+SS80
yvrt7RJJXqQ0EL/fdPl5mRnzWBLZ3Zkh633EVzr4tlZ3/7gCyaKYPAGeeEnc6I+jm+5n4r/Os3DJ
zzTEUaBUNideMyC1kSpSSXibitCUpOeSaIDUoOEm2Y0dTitwTnh14MKfD6zPYmBL3rrHXmqtI9Su
Xw1LkC53tNoZTtZm+NgKHcD4E6QnLErLX8eIddRwgzb/mIx8VNzEL9JV/HPwcfQKsXXzqWvXk88E
bGBQN+eZlGkgrVjpL6FINF/MJ4ANAZXuXDWqa4i3bnTirP/4Qk40pYgiurDmhHovl+V2F8lN0NFZ
j7+A+cZr4n8O+deYZA0JkfMKQZeNRCzT7Cs0XIyR5+xoM0TH5HAsZH8oJ5KAxgahprdyaqU1GZj6
E5//ujsdz4nfK6rSAbiqwbImPVmkLwhVWO9DAElX5TPL/Um8HI9n5xHNB9hJoAXPYx4QcqSNm399
Htf8WgHxL0JPoIgjzBcZABx/p8rV7/HYdbQj1tCgAgXQhNk4AER+JXRpDIENwwu3NMqIErxH3qzl
LWA9toYz63KZGcSmB07FQCPQE+F4esahbPZtcuXxtcFqcvgRs1+9SJufgwFGahZcQoqIVkN6YSMZ
HJOJD+B3y+7Id9SQY+5XbZ3lX6IIJTqbeZAAmvB3FmHzI6DUMh3QFK7Mdn1FBVhMTquwoluMrZlo
85BRxftJQJ3AUm64vMcn4mVAfGIwmQxUgyx5awisJ1uR5hDZ9psBQgODD6pjghMc4iHE5u14I2D2
PGurM1eayJBz0FG0BZoKQxioZLyRLn3n8hnKJCXYQTtHXT/ZHcybxNyCuRWJhRkgm4p07IWlQ+yX
+zttsBtx6Ps7EUBDbYrtpAPUSqgro1XmGe9A7UBozWSyjhbgPmH1tvCocBEgPir5X8jBQqbDxQQ8
7Wiq+aPx6ljZiSzvjmdf6m1xZLNM3vUaPnUf9OlITlsVfZivGCzxeg/vxuiVneIXM9wVC1PvLJPo
m6WO2yh5t59brvTHhPJZtlQBg79fkkEPQm6oW35upb0T5d7efmVHGwX0NZ+vPkRtxTUSGhXWuBJz
gjm7QRfmaYvvLEEb3QkYOhvtShNvaP8Dx/s3pJANd/rEzpQiuqoVwVnBBe4T3vIhC0ClPQHJx0Rg
ckeriuSiNivG7tE5nbmXGoIresXXEmyacY1UnvDP6eSVanz932H4Daov3VoSeNY8LxSrcbq7C+cx
Lz1fDnfZDh0CyMK2ORsFNy8EIpVLmmr1EVLaysxPwXL2mujx689wvf15LyQEC17z6m0tHg2c8YaD
cZQ9Zb2ElVSTeAq7ZCcH8MOFLyOoWcCeVN1BvRThKOI0K8jfDcoAkpyvxbN7U/RXRPqfb+s+34JF
8zelrbywGh9Sri5t949zQz1ysoNSMNsWD9G23V1qrmia3m5qXHVAIEvHMu0Xafc3U9hP99uIMCz3
N1ygh6fErYm1EZox6Y+4nNdidc8fjz2SU9wlDcNC1xpr+M22eAzlHpd7POrXFOuNQlV2FRz8ALYc
fSooja4CP8eXpv0lN0PVU9ICU/KUn6sc4CJ9s7xb2Ab0Gh+ntKFmq9sb7xlSaxzhuuIR81oZaGlZ
amvHv4YxYZ+d2Ialfd8+dtDKz+kUYG95a6rQf1ZrZpkzF62gtcGfNUsSFvhkulVDTOsmU/ZQIRUp
N3MLVlk6nY/t3O8YPRhjM+6wRSc+9SJXfYw3OSD4/zzNMuHlNMg9HieCKcIug9+NT+k5QzHLS2AI
CrpUo0wozqghVS6dyQXW9m7R9Ah/JCMuxz0y6Ybw8jZRXq4mDlska18HGhjqg8ZQ6BWcUGA8y1Hy
Am6J5V1mwhmTvjay24lGBDHjjKV46Uh6A9fk4oqLU5DsLROOSYHE0HlFtmJCZAptwHl21T3gpQGe
AykN01mMt7iZYh3DIrufDz5IkuQfREKRw2B7sTaswK3UE3BiakgZ/5D5El7qa4WspPQ4Njp0moKC
bp28ybNlmmEuFiEaHgm5/UpDfYtetdh48SLRwwViLINWzSIMLD6kKozENANimkkTCVk9SlJ9WSHX
HNxC7H6KVii4/3Ywi+YnyvgW6W71SEYYzHUEXL0JiWnvlSKt5Ydz0gKw2OdRtC6dvuvDyCzQnQi1
MgaiS0CCm0OPUmkTKCWSpFj3t2qbWB5TDKDx4IocdfGKVm5SQ2otoMamSBDWYYoDFwnZEUjp+xWi
gYCoSxx5k1XcMqzs4jFDXh8xNEHC7m7BQliDzsTIx188yED50T76qm79DBPUKzCTo6+sA544/ynR
2zsB3VkGjYdut896lyQ8EenjYJcfbebgCdu1s1SwM7m59RJdYuUO6v9H7ckKCgF+fQ5knWSqe0x+
YNZLkeax1DbDE7ERw5s6rcokeZpofjNujRuMjbwPM/I49oRypw/DrgeVO1229A4yMXXiH8QhOkaF
SsSUfi328JtJIF0Byk2MzrR09eW+9osX1aXLoyySCM+QjlS5iPtrFFqGv8ZxEUh3swjUQHpc/jiu
18Ec9Cs68XmQ/uDued7Gr+bhopHqvkWDzUkHp7fzwfyR523Lp13V2jtKdGGhCrKDcXEPbJlGroHA
gAJObkqbjB3cTozkOB25E6Zya+vjI9Hn/a96uhzGRNT4jUCshNq5XJ8inJocXwqAx5O1B/V/njpT
mCBrd2M8nuxmFYpaMw536ioemYcUc02enkdJ+aAGYd5WKkktQtuyDs4ViATUu6oSowgZI8m0FpCq
2ZCvjftUG231lBesphvEkEEB7kAf2xPh6/+bCGx6yp4lGURxLvEazlRIA4Qzc5ezRne9fWFX84z7
M98TyUYccs0+YqjLRXlSNIJID/F7YUB5adZmpB4T9UyRdfP/5onaTBVN/vMJHFcv4WAPa5sqVntT
ZX1ygbCmQxEU0oFKr48zjEsIXNiOi8ByIEzVrUd/bbu5bxTBsovPZKtrjCtyDFLdXRV7z5g8+XVO
ScyZU2nETqumUAl5KQUCytVEyEmoB3L0+SHXu6ftHnZLS5LfTtJ6BYm47THz2zZXWiqRP4H9hEGW
RljCj9Bgbmtlw1tCgPn2loItg4PZCo/e8WajPugebJvH2x+x5tZLRWHytQ07e5snvDJ8PNlkqy4T
N4IYpUNHI7tiLAlXt8b1TBVZFVrSUs/R67UBhSMmEsTe7BVo1Zo3DxEXNU2uAjNfVXvGi67heOaa
o2mHYrJnrv4N6+nM8BCftntxmF4249+g6Qo0qUC5fY/IS/I06RHu8TkvXgaz9W7NQHL4H2SLsrxP
poGYiWfkXCVkhbDzXYX+FYUTHznmkAln4x1UQYYTgD8JgPqKYerBISDRGE575f937hPFzttX6yct
ca8hQWlbpFLRott8VvNOlt6nuL6PJVIRJxgJe9y4FH4lQGXAuXs+GY6UBy25D5ltMY43pApCYZAi
8xc4XMWGyAc1q4OkDb6Z8f1LflcMj2tTksOJm4U89U49oNwhs+SiVAU4lllJ5LTN7u1msgl1WkgX
fYQ994BG0CrjGLg2XTMcRqHNDOYrFzvzb3sSFO9C5P3ByGiIowxlfUpFS780bzjOhR4r2yLHLD7F
HO+mh6TOaJTmcPeIXF0kX3iXYOXVZscZNE9hMj+eDIzAnQ6gGYULWA+PXocf4B9eK8IJZKA0AQ9M
M1QPp7O9EBWhrY9rYMwECvxUkOsudmYfuN06bARAkQP2mF6uAbj6cp3GZC50G2em0n5pzf0uPO+G
mCzZj4ToqRmFXgIWJUxAG2h7B6ZkULh4/k9t6Z6oVVMskw4yaobJa4PQ8Eb9ZPEZeTOW+7lgWVRi
UO6W9Yj4qzDQ30r2vOoEhN3TUsteBDmcsFm0goz0MJxo+1sExmkwQRXg8seRpdBcWzGxGAuG0r3a
bvL4Y81nkEtgzqUSsBLfaQZq0zKuEvwUe+79Nod1uC+tVa+5sczQJLRAwrcRanHwhWeHWiRjdU49
r81pefxz1l4fhazYbQ6W1QVhCNq3IlMttMdEqXxnzWNtLAeRQbS+uY4Z36bGSpesxak/fG8rtom3
0wheSYNpoYMFtRUmCNc2sArOIdorHUhAmLaz7T2GKc7y83sFMgYi/JvYnz5fNjzRaHX0uYfBImjv
na/19HFk9i/VyqLunWR7SLf5jwQtRg/VS9NNjJ/uYMdJxYu5jYXkwJosjYrkKsBcY17V00mEZhk9
5wEbR/U6+qmMeUF3X1ouqgbSrAFTNBZIyOU962q3L8CUhkLimacmffSVOI5bPOofOGD1iToTUtjF
vAVuiv9rJXoL+POv9UGyR6qZ7t9CP6JVSsZXOtyLWHf63Bke2Vmke9lQV1UkxrjnXhc3h5mTd1Av
7Djjg5LTkogmUUYkh+7Raknc8iMcruE/HWe2OG8V+01XiNcLUGYTS0kQ7kVQiCLevQ+le+5fbjHf
x5yTszgdQ4B/xdt1AAZyJ42PBicfYefbZgK5avkJmNv/g9sdFAspkKHaSSaQj6hkPCkaADOPDH1N
8SZE7DlKiX/3nFDj8pNrOmVH20nxdTF7xyw3brsMjNXdFgfZkR+1koSxdoMFYf8OfaJYj/+gBxl5
Gf3Xe+CdLqQ3n3QU4rVlpwa99CuCyyDbRpbS8h2kLUm1M5CLhXDOZxQH1eqD64VLLEXi3V+xWk9Z
k+c108fwoAf7DsjQEzriyyInxbTEFzi+U2j0u0Lm11Fj69s8knbqcy7jeALDsv67e1NdGDsQ+p9v
DDO06YP+IXeVeMNCl73u41HFSsmtGhWXVz1BYqWm3pT3l0watCOWsOpjOR3Ymw2pFSLbVhqZEgE+
geW4TgiBDtfJB8qjHUuB03RFWhd/ru5jODh9htOjCVX5pkbEyaMU9xlBk5FfJvcCL9TIyDwSE5xr
HOVwdyNYQctch98INiArVRKCgUtm0AxeusssUsrey9oVLS8EMhiui+cAZE6UxHrEW20iMVnwBUWc
OsEw5bjHxDV3D60CDyu3HvDAYp7W/u3iy/UoHPt7PVy5JyjybmIf8Aw5lFx4KczL5ifasoLLOjK/
x/8a4DUgtVt4+GS0Du82gNStTgrPSIvs4LXOcKa6UMonA/VuDh+g9MAceHjzliJHxh+UiM3L9IAx
stb7PfTHiIFgA0Od2907Mv66JmKyVtoUKAe/w78KJnkV80KznjazDzmXnkWpDk0lVvHkDGRhq1dD
QoPIxA+NhC2sEOkjGnpFV0gdn2k9nB4FU1muNvoFMe/J4JFKrlzeuLvWJ7A8hRmaR0G6+8W93ZfH
5HLm2c7EO9xey9M54UEgDLz4P+hAHDz+dheAeRcjuFR53NpA9DBPZszHkkQ8o3rtQiuaXgZK0Ipe
e+IPve17lK5WMB2gSl1v6WtOsFJMrLi6kMIhNl36WsfjWyNBkmqMzk1aGHaFZeb5e0T9Y6yKYmN4
KH034wvdhsEysVxlpo+sE5tJvsaaYwxvd9fnibG9sAsfJ3ZrIdaEz0dxfiTupVRV65inNbf/tU3O
SvoKrOuVcbHYPomsB/a5MOCGGY4k9Lys1hO2SCp1vEyZo9Yb7338Z2JqKs0VsLvjSmGTOgllKvZe
6Y0tt+yNE38jnYyLXhUXozjWkx4xvSzu+zm5qjw+hycJJEJNtm7/FQL9Tqv9OpC3Bq6k1jsYVPw4
ise4n+rLLoPtx9RLd5RRcMpIUpivEYea25l5K8UfPV6YXyX1ki2/+r8a+NSJFwefztf61pAlVAlw
haoJjUTcz9jQmhpv/BAM4M+nG0+PGptBAenmohS/MLlwQlqgzBqBn5r8RLu+yAjpopCNfou6e3Gp
/1SPOP6PUfyD88l2WRhkmH6VwPyMrGOIeBp+fwa6rXjdTs2N/PjA2bnTsNL8GMIDwofSZDbalv+N
/WgK4tL2odxP57BiBu5dx1BMcdmehpBEz1hi9I4lfzjmKGaPEGj4EXBkK4vkyVDxOyoLv7TIovFx
niCocOEA4Gp9YjSIXZ7eb0BeIJNZa8JrvaPriHU9xbpAn/Dg+Fq3jIwsopP+LbzGmg+eQq1QuxvF
WiAkswvgnRtFFRxtMfWvWDdAJM3C4O+9pw/ya6UfZ3uqfCgX3sgZp7bRlrht5i5nn+90wuZoTa87
F2xyxGi9yklzrBGvfTsWb4JLljhk+zlfmlRkWmUhkpSl94oxoxWNKkTxnhyT4hem/tpYT2GQYweK
u6oDz/abtRTfffHb+sFKwXIqg0XTd7eVIuYhAO25u0u2XPp2Quq8wRT9sXaxyLTZHR2FnIIlplop
1hyCSEG2CeS77e6jmtC5dvbfULO2596FItKfyMhp2vbOlMRjp1RZKNH/a/zyvQsycp8GI+IOl9PX
HRdAo8JVzMPSOHVzHthH4HZhc64z3JzP6R6d8d+t71VpoJr1hC1uZT27dy0GOwL7ziakoEY1TExE
7tsbI4MukYhxJr0IBTDZtg0tF8pNW3ilunpDhVvQGySrzL6id5tcq8AS6lHokgiEVzCdAyzGanN5
uUD8XBK98XOwj0c9pXZc39Ta4/T4m2p7oqRr9HFFA7R5JPNYeWOaRlh74BXe9j9WmLYxBmnzddWl
+zlfCMd4tPYAF2SHe+B8d5l4bmuv0G9fv3pnXKCIXTqB9wpD1UiLXjCu0Lyjf/4rsScwbdkctkPv
tWWLC/CBv9tVGttREW95A92MW7Wm01W09Evx51u8mijbcqgu7/m2wE+eUyML0jSAWdkNXUBB6jZW
E55/RxtdzZZ4O29lQetl5G/uW63vL0f8WvXc/zJShDTi3AZI5yFNxjFE0L+awo3NEmjb3Jh0nFlY
8ljg71a0OK18Ot8EBVgAkycB5oa8WrNv0PxMkr1RG78piN0mdW7S83Qn7pU3mcXCQ1y4zKHcw3z1
lZKRiPoTvfjPlAArSFtRrRJxCYO4pKYuZi0ZMfywZgWC4XmUzhsgKOy1g9vf1BOsKQWcrUzxMMn5
gQkhYvpTAT8wvgdUmYMETOJAym/WjLeNLfamSvFR4m72k7lQvvdLhJrcn9gyaziq5pcmit0YtAuJ
QBxV8wFsTcBxtqzXwlKn5TSHbiRVSecAykhvU5koST3vsVWqy4d0T9tHTVqMIJ3OBqkW3bchLEDB
vSSBI1FGMeN0Vplefbswrmm6qtvoSHg1YVKLkJlPzqK/xGMPQt3wsHgV3lD8FnwUpirYyBRAhkG2
r1pZH2oMWYr0i/VF9lbPUxLTHOIZF9QQKzJGWkffGqzdTMh7TyAHgMF8nWfvyJjlDt5kYQfp1gLP
UXUt3urfUKhNl2Pc1RRtq1A/thPaaAb3WzN6crvQ1ZAxvePNjgZtOPuU+i8r0jta/he+YW24yrhl
YLWn0tyr5ymNTMJ2P8B7MdoKjxvcy9xqArd7LsOVhOW0dBu/zKAIvpMslwKJsdKvDSaI72+qNqU6
LyNE8GXTt54adlVFvnk9YdZ5luG1q8JJGlpuxOwipf4F1VuuJf07Pw5If3hJ4kEqtaNh2zuhXALY
nd94sbayBrPsJbKLzfEu53yjk9OEbuybSYT6Hx7lwqdbx46va0Jl8JoKdquZcjxO8xThoozBcdpn
GJLc940Zsxlt8FOemuOKuN2gbi0Z6wZkOZXnYKdd7KooNONUBs7Wd+5MeRWG37LzmvWPoyvYF9iU
BFo/EalP7aTWux7wgCwYu+/qQIyA9kfDVVKzSPXUkwsqhNjVbJ+CKNDBUpTV8pkSMxqRfDYrySM+
8mgPSKXz1RLpHQl50OUczWO11q9iqpkdnj/t61MwR9gE95UZPrOUMTtvm6sydH7eMM7aoKRSQKnY
6dXLOzUoN8T07iizqaDWFSUWYcgCoLiULRdu+t5+ECgCCkiJat4KhiKlejCntWvCxSAUhqVqBIvJ
2y7Zew+P76JuJkR8FnBZjtfcd+rW6UgyncEcU55ClzyOAhMnYi67oVirq0d0HTWtuKYo2lvFf0wa
/sO9bfXmyg36UUwhTTU7xTAvM0D5QFYYrZRKGSOZO/KdFofw8ZYKPuCYSzrZHJR5O5zsQPvNvlXW
gpEcdo9EcWzOWMYZuc1N5aF6gDCC+/8rEgjwy3E328TysHLjhOUSUDUMJhuRAdx6N1rZORLP9Nub
NIOmCSqjQhfImPukJ7iYYcSU1LYVLx5FA42M+Pv116UPLk8Rccg8KOHOzgbsGJHvzS2YgpZDiDlF
XsI01wHCD8OxSmmGxkPUjWxBsmXtLezlY4osLIMGI89MBkvK1HXKqW4QiYWgFguEnaSsCH23w8k2
cj2KiQtgbPOVuhmWm7suV8fOG73OgB8CZoZ7U772CrsWu4DDKCAbc8+JKTm3H8gQr9tWQANRpd4z
x2KEvSNUutiP4cTnCOoVgoH/yFegzu+fwsAqu4ei3hbn65E1ih13ssXhhwBP7HWbkpM6uVBdUuFp
hIVaild3ZbyDIb7VRuV9OSeL/0vQc2wXRoRFLsnrsmQvvODVO+mz36fOzw/e7zvqiETYtBnS6wSV
CA4GUtSpIsAJlM9hKITGq7VkBhHxQt6eZBGNva6sBHhIpzHMyQYktFu6jCaOveatNJaW7X96gzyJ
6YFqEwbrvKmRF57hGljRikMOiXvLWhqu0N5gGf7Y3yJ3Ka9YpX/7Id7PHswDVmkxA8SCUNQHVQdr
wa70WkYJytlyzaUEUafkbxuNNOUJaVpph37A6MIIm4yp4WuVK0aveLA7eXVNELG7hYQAQewLEKyf
h1rSJ5gGpDdvq5JIZSMH3bvtgr0LeS6++/cgvF1jeh0l85Je9qdzNWpesvyca/V10TankVM3vLSL
krrvXlz0E3eMj4DbKioKsrwkJ9QlKw3Fag329TY/MV98hbv68KdYP+Sm5LNwePrZOICTayTbKxuj
a3WQ7jj/h1UAYjU52u6KNX1ZnSvxzYkzY037dZQRt6+ckdKNLfcWWQVZylq37X+doaHg7ZuoJYw5
3FAGDfl8zD8ytABCWZe6OB+aGSsTQSvR0j9wsFldzwFv0xIz+rmACVSXdTfIZXNiXAVafrf3vuLJ
nV2Eu3w8YOd0yJd7Z1ELh9Aqd/+IKaojgjje5+ySXZg/Hmpe6deBRK0M1D1mkq2NNZ3mfZkLgH4g
zhr/nzYCZBP8Qqsv+l85I5caO9fTIGiWZ88SnMJWW7J0yUFuI6/9V++C0n/F+Fd+ICL5j5NzSI5C
J1lK6yILRndvh3w89K2hyo9FD2nyVmPN0rF8+cbdWG7xrFWDBiWw/W4eIPWB54cH/BpU9UIIDll0
ZYagbp+LsQejw+76gnnoc851/dbApfU5L4rvX4B9hZ9TV4trymCE0JhB1M5JA6hCZeLFLO5BaX5o
r1AmW1h5AUT+JDx1Cs8KoRVoxVWnnMTPkasorTnWhBWpVW/QP5rmfP95Ui+BT+W0I2y5RQT76mdd
Rob5pQk025ZD6aTKg5ag1QwEQguOKJdR4ErHMFc3B3U7L8clvVn0nhy9e+NjLtdE4DQ2t4ZDVNIi
Yj0BrZREmScbBj8jwvOWzaJKeeRRjuFhHWY7QAmMGtv/YlBZRRe67V/jKp1atuo8GHQ1PzBG4ihC
4XYVoDEGdgs5Z+0ieRa8UudhuJmBFiTs5R6lmqgy71qBdO5TzlCMT1TF9SREpcKdOno1cePLUe01
MAGKSJBiKTSmsrCRE7zKxhXRB8bV1YZv1hGOKrv1syaIkyTxdeV3a2H8de8IKt/vjc5Zdh85N484
bDM/Yx917HTDqGq7WsfLkrZx50C0U8W56aE/Wdv0borkZDsjr3P8ko2LZEPJvOFB5GWqmzyw6cdE
ZNwNMtci6sDpxCO4VVGT+DVvBbIombOl/1RBJ+HQNhOY0Ih5Qj6PaQ1TQGe88q5bF/9LBW5AWjKE
Rh1ado7GEUEP9ss8nVlqc8J6+Ev3oRhZ9qHfVuU45tUmoOUUxZ1IxfJZ0YN1kK2TtPF0RzD12LNE
7m/IozR5IK0BGDAbiRB8XDOwsWJMJf6iL3leLlFhXCvd4aY5ktLpYYsu68ZSKWBa0ayLjTL9nWoY
wsZquPgAR89ShM7JFF2I78Ng+VSh58qu8q9PtBGJek2y2RZc35fjlJl51x9TujLf7Cvj9eFFDfpl
hzcDSmfdQSbg3gmAzG8Jyaoj3BKZk3gu/CPCzlqV+oXvaRhcdWCjWZEcYGqJdQLSisziBPLpHvqG
Yunoga3TnnQlQkw/ggIx6XiiS/y6UQbPKzFEiZ2X9Y2tc+sTGPcNwJRwoalEroruvR2gCyiWE2xq
Qasw/VkCA+PjOpnVfNFtwFKKhEIfrWvEM0Hetj4gqLCWELbH95QgCw1Sqjgol5uZZtxK20oM8bgu
Kp/v2h0BiSTheI3UE0WzyXoQKhgrGTI6ftiyVwoFqumaFMsj7Kt1ymHW40K/5oJxicRLyyxDgRPH
QX8jIdim0F7Q1BzGty3V/0ZXIqhhz5MiWh26XIE1p6I2nvRRo6ERYU4IR2znPGugzIHMnjf6hHtv
QWlxk+oDyZ8UXQLOfeDZPLO20OMFJcZ5SBpYPNhHeH9BK7B1MUkOyTXy9968j2e/xwGwPrQbnB/a
Vs6YMP38SSyNEg0inyD5wUJDWtP+2v4GC3WpN3VLqgPJOH8hJSO95aKC3asMwJ0Zi8y3iQ++dWtx
da2nT1Q30PApBZbIkjGD3t8FuAtLEnBFwt0TtnyNT9IChHVfk0TfagAS7WVSmhea825HpUoYjPhp
xu7BjmZnXg75jrurCwj8i+PTavPZ6IrlmUFlDWi3QORLX8GQdrsfxIEmHC5MCmTUDOc9Iv0w3Vdt
byEoFFZOcaDyQupIGJszGG8yiP55I0UZRpI2lpOTJwg8gvv4j/WQLh5lMeNm+6UyrDa3d1TLvZyy
Nk9FphCPp4a180YWnZ4o+C+wz0R6RAbHbWm/vhhObzQyxKeCv9ZjtuEJKCPSvINTI2BgZzFCtxwo
66u1Iu40AFLzmrMc9LalR72lpNhRi9Y41q6DoEOf9jRSro5E+jKNOdrICcx2Kz4PYpiEL3YUjSZ5
Ul0aP5qcJXhDT0Ojr8Ksbxn0gctdPbOwwCYFNR2GNo/1eUk2qiX3MgaR8g1fTJIow7w9cYl9aSlV
JClsPYppJGzhfWHfbyq4mWYYPBvsZzoM7A9vwNllMSUCHu3DpIT+YMvLV3dHKQpf+Ar9yAMm+bE7
ERL0SuqPac/JSnX6tTo+QRjBPdsrasUIJCrXzFPBolNjjgg9mDPhrZ4zYfUA7yje544Y83zNpffc
clR0tiN3OoQrpY4ls8auGvjYyV7LT39YtQK1FvfnjLYaGHFp1JW8HPtQRCR6iJwHCP5ihS3evbsc
J7huWwm6V8wAV6bIrmN90MPXTJ6m1Ac3SrBx/y1akmsVMvGwacNhRXPpUo1mG57N5fwed7fWzNM+
h4PO6o9J7NfX8GkVmpPz8uSIRXUR19+y+gXw70oDaPTiv9I1mzaOagbN/jN4SsaAG0ArEKPvCO8m
tNOE45fjxabKMcxfXPyQ3W3kBBzuGGW6BYg+7NVQUb841kWdDFQ8EAT6wsxTsm8/EjYZxfXNt0wv
lM67Xv6Rvvbaem6lpntPJNYuC+d9hYXZHnXCRnNcQqtBOWJH6iMioMDO0t+Uc1DrWTBonhbg4JTG
w/CRHwNtHFMJ7ZzNfakFaVhiEo/hg2O7lcAPWCedqUFu28FtUIfsZ/0kwGzHvDQY+vGN+qc9dGzN
fRs60DVP6ViXnvZr+V5buEwPrYWTBk/Y1rg1xstKCCW+t/wnuKpOrWomIaCzZ6EEQ9x4zj/xrcHb
oJpfKvDL0gppYW/09AxALwfzazjzW/VhQMLrAIaKeBD59lCTCE3zqKJf5TbUCMxtUvBg2chI/hu1
Enhx0iBx8qdZJBbzjzVOMDiBBO/cI3GyEOeh9NQ7PwkKQxyi+TEN/N5Tvbda1ixhbWJbo6jS3FL8
iHcugqzDewQ8vLileL1cpIdh5Et4uWVEBaol84jiKQt1ka5oujOVjXT6EOlBxBQcXE9MPmsSEoMQ
3DZyzMFu6VmgwVihlwf9nBm28ZhO8lfXTaxObbgbopnA4Ej482sH0o140VGugU8q3iLVS2ipa5nx
CzosuWL3/fFCuCFISp2bQzXJFkrVwWyCk2pM9e+ZhI6oXQUJE+GM9rMdp3GtarldvDJPSNvtmX03
LyU4pYfAZ860mc89Kn3UYCfpJ8M/vUi/l4FpceMLMO+otm/7H13Nfe15MuaYaUDhrTnDa6uLI3Fy
w/4pXXtcmpNIZVJsyGiBe8TgKef5U0QW0N6QwKixXze6yPBv3BdctR9uqlogLsgOnI3vBoNjDBPi
WwKBpqIj3fmUD0qU1qCTgixzEn06dzrWsQAoayvfjVM1qLacJDN6fDYzldGS0s2nJa/gm0rndz8o
dW8sKnmfuXgLcwO/FS0pdyTIHXMjGlaziLs9UcoPCYwoyA6jD+SRZMynQNX93nUa7AM/WXpOZ6RQ
YT4dnSefnAPcvqkzkaWph4q2ynkxtq7hjuNUO+jsK1u/DRXYDdgbA0zwJR9UTT3XLr848BIknJmQ
ZjHN2kDik3I/LX8PUzh7HDkw4ENYRP5jvIZydnxhlGZuKQY/uEmA2XDfDgyoFkPAihOEW1hsNuED
H9tqVx5OwQ1/XFICsWe1X/0cmWy3S4ES9sOGncZa0ZVn/Oa5ZJeMMLqwWeaNXMaXseMtsygtpMWM
PrBoB4AsB+NGnGi0SWkHlFiy622umf7qHjVtZpzgZKA8zyixhSi7JY/PiWWlCO02D+E4+49/dMSh
G/bfII4VZJ/ceZZmAebI4TURHBX+BK9MgrwEiy41nmdaBg3wtoXxrwnMzo4w30Oc0E8L0PyPgFJT
Bg/LAch3/RO3EwWyife29tNB+e/sGoU3OqewtGKHGT8Ligt6A/1nfV52SvqtVispWao/EzHGB81E
xguI2InBy23rExOO8i/fVKldd7A9W/yMsJYHMavsDNra5mA7lvdwnjF+vZiNW42PpSdCSbqf5g+P
Le4w0eSzqYY43ydYPHmkajx0JxQoJB6HicxpoSrEo5TR1RB923oRFSBtjVeKl0kUEW7l0ooL1DIg
9O3RNEE9ei0XWzeNoBdkMiT8MpUJa1TAY4yKbezYjJFNzMUCQ4rkDV2bOij16OW1HhQquOHAAeem
Kw8hK9HNJBwEWEUYcyF9iqJHU6O8ypX1R390bEPNlL6KDSHwaQfTfgTl74FlIu9BH0H4TII4RigI
xniOtC94eYQ/LnwZDWaf5ecgP6aVpcYn3erjjo0x9IJVU+Ndv5pgFn0yUu8lAK/ypBcADTGuzv6W
f75rpoWFBW11jZmztSY3GyciuzD3IxXFV2M4hoGjX0XfXzIJeYkPh3jxBOo7AjHOc7kqgHKc3Qg7
6FJIYxb5I6Z1Mtu+7ebwrvsE28mwMl1lfmfjiznJFDFrMMQh3RrL6nyajcdfWtWqGt4GAOYGeXim
2lyLBAtJoqGlnftDSMJRLeDBA3u9NLRhuVA+2tsOlJZWftx881wVSEq+VKS5bFoUpEFOKvh76mwJ
dcIeH/tTXup07mk9oPCGVmdhfObmdY0UYbm0HnIrDFcatBakfwtbeNNciS8NAGD5zVm0ZC7uUstk
xthiJVARdwU9fNNYpL1bauakY++KAGO1eq2h2AptkYJRlDMQdVA5+hyvN1RBB5ZfOvwACC7juELu
Xm3o7bnKjFq+Ye9cpXWEJ46iptPl1QCZTF778BCazLM60x7WR6qWCvfEJBQLYBxyKI6UfbuSvRwc
duSXkbneYDzsAvhRhpnLb1pc4jOq97trN1beTj0btxhyPmScvD94jkrp05MtAOThYX9S/eH9k6Ld
Y8IGiVl96vsaaRmOWPWZxQQmNaak/GRzeuQSIeimYkdHL4/Lq1I2/R9kttEKZJKpn/H7pSm68JL9
pCZ4KiB2XJ3lFV5jfDNLvcROVdyADamFVm8lOY96PNhMoc8Ig/9VEf5M3nhHldOhiWxjqiwT/46D
aYo7zSmxYUO5IJtzegvwzie6ywygMvYMpzm1PocyVAo+T+ekp/NtuxI8JukF8Lnxl4nmL07dznGl
zsuytM8XhH7rbxrrwe2dxnyY15qNe/nK39U/HUtVKluYVew4gCTM/jdy6Rpkim2m1PgJilHdV+t4
UaV9Ul5YaLIt6yo4OC6+zBYXLVFxiUP0a7a4uH+YHrY69NPCDK/OgHMwB5pLsMJQlfFfZlf9oCSm
X6OjMQsc+IpzcT1dOcaR0CwU4zRgOUQ8ng3FDh959+Mz9a/aHpyggFn0v+qw0pnyvBwlMwS8IMDh
+T5QkEFidyd/IyXyLlhRxPMzqvJKl5rnuGjS0xB3uFvMpE3OnxMtH8NM3GYbTR3rVcbq3+yH34Sb
h0E75x0sv3K9zUmfhkqhae5+foFOtuRAPE2LO2jBjNet5RhR3ffMqtjOAdZX12h1/zZI6HwSucAT
/RAwT73u04mrbOkp2rzQYy8305liIXh6lhNqKSWAO/clnQnySph+aY9E2MkF99mTeVuDaKK3QXaW
UIvRz2c3kQyPb2xNOWf3h3nZMKI7hq1WBu1qgAzgV7K0+8RQs0f9YYHkzzWJ6fz2i7714zjoxNB7
ZA+HnCpGjx5vWBKKRtzGeJ9FuLL496i6xXIuC6bZfSJLEjQYMq4Rda50pKVNHNHvYWHBGWNouG9u
FeM3OuKQLVJtmX60XwWTSAOjZgKRz570Gotaainlr0Rp3595LMLcM/b9kWKnrFiduv1k/rdILBSZ
Ut+AMcwG+tevJ3FmKt5mnUa8enuWxNEfKt2UJnS4F3ahU/xPQa0/z8vV0KGUQHs3/xvwxTEpQVMC
evyn4PEXgahElVMAFu3JrF47NY8KHddtSZP8mVlI4KwyheHCaDu6EhvKLNoUvmCzZ7P0vCQT9s+2
0ONjs/n8V+HDC7Tb6/+NxqHEI+et+Kbv46EvfuZCU+fX5cK08p2xi78elJVWSNgeauLOjxxdxiR1
WQkXRHZUy2ez0uIEvoZf/0G6PCZdJQIrU67TpfOK+NOr48YiavWxCKluJ6w8YEeaNzjbQa+QvoYo
f6vVmOkxaznjd6KP+KFej5q4N94VIT9Nd49bulDtLtTtSIMrl48fTOJzfzWSiYA3NULY57wSita9
K2Znhtu305f/qvq3QJOv24TpHR8HAm43ehYZgQpjvC0lm+eYz4N6IslO9hG0fVp5GnhJyuzaBAZk
8x/FLqkJm82pUlEcKLkn8Esmj8Q0690/cpUZQh0TttrWmAzR+7Xydw688spNNI1H3opp37lqci9Y
N3tRvugWRcaXRtBfCj4+7lZjlw2LGfYDRPzc752yAPU5dTZeCrgLb4jwbi608OpQwKdOM4H/zDiH
7R5xs4ivguQ9MCyM6CPqHCvlDCWxaUWzd68qy6oXn4QJsUvzScbewxIx9pBQg56YbZh3FAZ/9vGr
fphTYhDQzH9c0ZHy0WWSXLnUC7EdAcH1s7j0RcXmM00UeTEnwED1nwL70fD1wHeulsIj0gW7Pn3c
iPGT4/ORUB/qmiIfu56EX2W9PR802uDP6vIS4NODFmWEvEG+addfQV9xMs+GWNmGJAQFJP7SiTsX
ZBcqeQjXGw+ecMQx/AzzKHyttsOGZnDcjh94GY4dsk9wnpx5ppBcgLXdIxHoqXp8mzNydYsAjRs7
wk3QrJYkXaPrC8BnXeRfEyROvqOFTAS5ePPw2OPPRD0Ts2di4zxUs34MGu+pKjL8q2cCgrpaM7KO
dxTYBDPgZM4lJxoxpxfjmbvt2grvW57mneXILgHIchlTewdNBPVMAmpsN5gfHVXE9qj6V+wvhczF
JGrcqFg3KdgcyKFHA1g518F6d+VOQBsiaERuAFHNaaF5GjO3+D1Kfm0NkEX6MPu9+vH9B5BA5AOU
aTHgcb77ZvXsTIak8iJM/Un7+PHkaMTMlqLDFnbeLEFq/wxh9AH6DQJoUaUD8EOCrNKO1rT8Icr8
UjD0JIc34K0PWj9Rd0aXAF4kg9rGZRhd+nnefZ0NMNDTNJweAuljAwttuKHYPBt/kOmZ+FyZk7EF
J0iYYmmcd1xbjsbh/Px2bXkOMG7slxuAjNOpTWoFhuUxqznf02h8FTYPUEhyKjoqxvxYQjvNGk8M
ZJhx+4vTDNIGQLkgr0ljK/IDMO4yk/K7PbmFzEEmslct1HpaMFCYzBESwJsjCRUt9cblTbKVDnHZ
WzuQvx7wFzYMor+zCp4rS2NWkyih41qvR335/C/rYxsqcF79wkrN/iGFZcwuDFy9rTXeWy1vFX2t
31TrqSmQDyU3sn4qLzGmf/oU2/l7/zusmU+8bcsyzYqbFPKIs1QgyiWAlt4Ne3aJyy4N70e3oSY5
9Fx/vsjS+uVoTSQsyguIOKT5uhRRkxW/TqHuPMxOgvAzgLNgKVYTDg8rxq5wIuO/hh5hFu7WTArA
OZN2GTxrQyXPoJ5U/oQvzoiI0QRZ7UUovUeK6nt7C5cXb9s6vu91wj8ohNsxVupEifMXTneTg8xc
CSQN5Ny/f4+i0Y4+O+7SiqDpPIrddkM9nfsKaiDsEAyfL4/adfY+8fytf70qsXvD7NiasUVbMEel
uojrTFmN/qtPanVmi1uvceg0Tmi2j+BLJnHstrFHWJzTJKbdXIpmgGnvPOabuExzRNIS9ahELp4m
CAd3cXw+/xQynRNfEAUAghmSe1Ib5Ee7qoPp7lzGPFJtOrpUGojgNzkB196BCcnSj58IPgQf6D7p
pZGjsFPn+2J4vZ4f4hbsLEfe4aG6M5LQHRBrBF+m79WANBefHl19LC/ii+DQMj6/Ikpm7KbKEVpw
o4JpW9m+x8Am37d6n538NtfBkzADUky8cigh4lmkV59u4uYYLTnzO0kO87YuoRJRMSzl72lGtY6+
4H1azoP7lYRAE2Ze3wqGAvjlrcOlqgXLm5uIdasoCuH0pPOl9avBZOu1FfMw2TOX/oFeYPxio0P7
m9Haz1xScDRnp7jbvwqCUGh5MKgy3zqHqCHXod0lLKBMRynDUeUdEzuY+zjJOj56KyURzQTnZ20H
Qx0N051UdfKW9HyOL2Zhs+6gu1G/6CFsqlSgmzhr9li+at49iGlLNtGdsdvhA4U8vfEmZoKrIXSA
hf8dmx1pHAn9ltjChsPQ7PlhzjI9gQOpzdL/g2NCmnmFhF8wy8qmb4S/79kBnaLu/DtgLiv8nztn
RXEup2kjlTo658hKN/KNpiBOdMAe5zgOwDqQVGTaWqt3CPoJ+7Th36Oy77aCpBp/xAbJAamNhcxg
0aIoWKuuvswK5Icm8lEeZ0X9EnIrESO0ji7h+h6+is4q7JW0XQ7fsPGIIj6ub1/yvZV89PWOzeSd
uKu6wsXtkpMHO+GT+Al5HXKO+cJw8afDs/ClATdaz15Q9Jd2jXMfj5+A6qDCXHMREdUwz5xnDBNg
skiXJYhlyi0PNzjN4Dom/jYfxxB7pi5qe8nLeLoxoV5v0KXbW2nvnuOVUNHDK0wHKks2HK3wzHug
7e2wlAHbw4lnx669v6qBjzvNy4WUOvWj6dQ+Q3kTT1yHhv+YenOs7214DKe9jJ6TwJR17XNp2eTl
Ug92P7yfqPwNv7lWiEzEp3ktQYPdG0YXNX55wiZ4dibPoNETzG9wtjEhHOB1aIZsavk2dOeM10iy
E5/N2oEO0yWIgVxUIgk/FcQ0cOSkcUj9V+2SP2b2uCrOPH5GB+VbP3naBnw8IRF0/JQudrAcq3hh
wXOXmToJkEapb0hndFm6lXE8gefKHLMqrQXkVkzeQf2uSnDiZcTC44MhbEjEry+nG5BLSH04QguF
IGP2a3fW9EEpgEu18CWz8B+GCYmSZW8OVmDONEItJUDB9V9gxWaT2dv+VP0ICLIJ3rdOxFx/IJbS
R4mUYJy5WRDaSvq4SgDq67afyaTvUC/jF0F5YSAu1jEHDqm/gaoYx6Lyshif7AmTm9EKDy8x3+vm
f54frlD+T8oPPbdQu5ua/Hs8jajFTd6DK1kEQNlAC4PnxAOdjIFvfl5H1ZnuUG8m9h9OzSsf6H1+
yGMs5uv0UVF821ZtxocJBmgNnOjwHKzbyX8Hs7w67iFTAi9fnF7E4QpkfNYLATpxP4S1eLLPEjuA
OZiWWjJ93dvxPa2Gr6V+eUvpeefJH/pkQtkluHij6vByirfDKfl3uQ1iNDtEbHjygBQiNrvQ+2zj
NdDZUNziccTQi41+/Wx5yU8ERB0fZ2zsPskzYCBxFRVcLjGemDh4y7sb6NllE/EbVUk6Y6TQ99qg
sTung869Nkmq27NcCfJ7d0MODX4xsVpmPsjDbs3XxOZ7z91kQZeOaXRBuU0Xs65u8WKvGI7kLG3z
Ib96Est7UIzJs3UigGtTdeD5U2AKGccbuUXSHU4+lxXZxzfPKzSSUZUrj1VbiH6kVVd/0s1PXxBt
2QIHnbt3aq4fh5TrC2TXdF/nhkVK1ThjQSUR1HUXWlLIZ8VUfUKmfMHRmV6EfFdPsiRA9nhhZ8BI
gCAp4m3qj44LQ0OTPwtbSIXlb815ggoHACO5Z3vUvWKswWezJsL1FNDTWWTn7G3+OtqCub5MJDAp
ASeDG40rNXTOPpvlI5wBcT7PPFVJST7UmW99qu17y+DvxQC1dF1yGOTQeQvbdblCNVmtIDGJpNCM
TVJoVR+pWo192U3YKf3lMPW/wuf5BfwbqOqPTzSAU7nxqHTVf3XUttefQP0JHStjURRgwv2CqMFB
T7YCOfYhWeek1ooMcRxEwM1rYPos7xkYs8QOA4p7sIPxS5KpCOBVQp+jiykFh25EL2t5/kEXm6Ru
pY1FPGVBVau1MlNHl1zbeg9+3xW1mbm+zMMR7TT1Qt8SzyeYXlcFrjUPMBHavdFuRAsyAkdyCwDh
o5Nez2lJq9ogsEY5UDL+EPuydu0p3Hthap979IhBsu1G8DLFZoRCjdYfVHFxBy4C4w/Tdgj/lHlg
syvfUqjjl01mESSY/Eh1AgCgynpWqD0Z1tWRqGQdzS5K0DvFIMEh3U8n3+4TflVhIe+Jsg/xbuLT
2QzQaJonEK7NZt10+tOmCcvw8Jw3emIw3AldtbPDnlJQLPwVu4XO+EuFervC8ZI5Tz7g/gOjRsDN
EJ0AQWaoeX8fsRYKZCpElaBNm5Q/0EM/xLm7ghkGM6ZNS8HOsGYq8bOA8HT2oiQQTaFVzk3bp8uG
fAaMk5lSo79TrNS2xjczNtvI6Z6SjW7UYiDVmeTElJPhMstHNhtjmnZv3slfZ28jnR4zFAPJxPHW
VmJF8nMF75dTolMVErWA1HaN+ZPSBPDQsCsSFBkCCgF5mUsdEiSCb9eiBOBZO1mFtA2pEsg8cRFf
XUT3IUwCoM2IsPQ1geFTEbvry+MXmKuW/RtB0cW2fvbtIP3Y6VHYAHL1Ibu+sazM5dVbFPIsQ6PB
7XLuKT1MsNzRBmRgbycq7m+IWC4FIjXsUjwXC5n5/FOOUCeZ3M+lPwpzXX6H3jqDqDY2RSecD/5Y
7Iu7XW8wIrkYAIucpKwwBPm7Zw1JRr75iTyb0Bwi699VgpVai+zZQodlVfsN+CI1MEDUTst3Fsc1
sTUTfRBBAQneSiLbEqsEvWLCOWHdcBtcF2CiF8qSshp2HOfA7flSsDFtbMlTp4VgjBaMyXpy/6QG
p/HEqjClzyEhXeF/VE4qWydp8L/n6+GI3Y2B1frMPY/x8HwcOC0Vf6HyCdbiiP28NfP6caf/I2wq
6kdWjbZMOJZ6nf9NTLQLtB7WY2ku9w6uvohSC9cVZv2SpOIlIdzQ9dzlsQPQ73JXJ+tpSl9uuiYg
qncBnF79Se+tfqlMIn0kqOLmaiLGWzAu40bw+fy2B242KcTh6ehKhH/Lw8AuESlWAxJnvfGTsmwW
TmBzs1mg0z6O2sRj23ra9b/eNqgyNMAKQn5EpkZOjvxS1pyF5LvYw0JVQuZqY1BbEiM4PSWfRyW8
DXjgucdKwS8OV1I9pp2RbVf056SYlfALOpsbUl4kvfKW3z0q4GCeIUFyXEuVOd3lGUf8vXxVY+Jd
Nvg84/EXPUO43iyA8e4aupm3jnPaDOdeeE7+RBJWHCLXsWd/U+/SSeo4kUXaKpbfkMzU9yRFb7QR
BxwrM0zcod/aPhNVgiIKRIzHS8zq+3vnVS6BmfReWVnBFMbySBq8/Fr71LQTXQbozSaHS2vOhh9h
f9/FZniT4nQD3dedbV7ugRRQ98i5iDovMwMvX/FXfWwsxZeBaihpcjZ2MCIwOmrcf9u4Dz8atjAO
avRmZjLApc2lTu/HsKZhlvReepS8GQRe4X22/687z1RqYZ1NEWQfdw/Miz2cAdf/sjpkUmtuu5Mp
GAlkne63YQnElWlwYUNcpUyZVBtbyC/XOJ0ycC6ewAXQ/a8beCGXia4K/1XhB98TTEPbzKl8B4T0
v8yvDuu6Xv/eqvxsl4QECUilgPSQRJVcVj+ilgqu+D+J0iUjVu0smhn9JfAalBv0FI0aAq2khB8Y
hBfiVE053pAnliA67SGySuEPitCTjHCzpl1mg1xVlwXhG/nSOJVRtP7n11vo8aY+vOAo1ajSCe+G
PVM9W27wIc0QAOaOxWlz6MS69QftkBaHdD28uiP3PGYMc/QKBjMfh8jF81iFrN6meOOTv2YEYgQx
6I250gYPSwy9ib+xQUjG6vz7pHNuKTIxLVoDnh1VVZrNA83fcXlV7UBjpzLugcbaBRybxwfXMP4t
6c0nSUGC0AY0UnB+KVo9v6Jm/cX0y6uQme1UCX9r47nwzhDtzRRPwbPQiQI1xHUFwgCoPzWNsOGH
4ioOuxcaAUGIc9Vec4+r06dWKU+mpzmlltXhdZm2O7JKXmyi2qqfEc3vlo6zAIRsFM8zD4v1iaQX
HxdX6imVdbTqXrDXeVa/KpV/xK7+zxa01PLGGJwbipvB+FvTddgFd5fKzUdEbxhusXtYmz0dDhFz
291unv3LScXHykbxsfzSUA1CD5d2KF12fUmI4Ef/JrWFNkZN7/S+SfuESQP/jaQ6ZjeWWt9CFrhC
z96SZQdx3Hg2OK5Lm3AePNy/2Xn1XDTcjk7v5zhAgGOHag6rtCJhqV6lxgplByIJOqpWE2CGeqbU
wpCvqhwtnRlHYzrpiXbtcjlGrqPxeq8cfJzoly7iJR+4zuGEsl4RkUZ4ptaetLfZTeEWt/uHAhI/
Icco2akChCmoQQ8ppARKwLP3hQw/tqyfKpa5/51RUtCBtxFSZajsRa2dwvIkEEQm0Zy75oS2pagz
5WUpKlWNFnlWGKoPeQ2Dpf/dvgSFOYaJlNNpA+GNKrMR53wkVdXBd4efAXXAnBLMCTrwV8Nel8Vg
LeCuu1gwLZDbMXz/ipU/a9JSMsluqF9aITLf9XKhHSP7aAK5HEj1aDcaKqSVL+KKPQ9wSa72zPKG
C3Y0jlLlkyiohGGBTi1xFaPQoYcdg2nS85fwxgdpN4GLlgqXE39YmxJgCSnRO8tnTqpuJUUDKKOM
OQ3YiXY+JEiuaVPIUJZbSQJHQzcOuuJ/BUeqWWWfFygu2D7tHV9xveNJWwf2rBz6S3NT8zmmzCsP
lC/iWZXH6OZR9J1Wp9YmKGJI4UUhDi1c2z30cvM4yL4Fc54eaY0/CW3vNi8ij8Avs+hmmhlWq1Zi
fYgIcMX0/rRz01RNSAwVZSLxKvvAZ2yowr0HtD3pVs9oq7oPbRbX2FyVPkYT7YOc4F41scWcv1wr
oJG4gMC0e7igLlVWqc05XRiPlw4Db8I4bdISLFN+vVdgSK7fYKl1QZnsOP37fPHdK5nhPoW3TQug
NfnNTx1XUD9vyTy0xMhI4lXlH8XVc11ztuzr1NOgsBAOXiMENYI5o0esnZVNXnfcQpaYLQZWNRNQ
Km8AK1tvIHBJ/wupuPSVXGUrw3dCJwy7HtD2goOwr36kE/xk40zLH3W6sHMuNeUiTX6BBglBkvb0
/Mfsvl7bkTOxLYhyIB2oBvvJv3BnSjy+5Fvn9PiXN5LwVPJXThdWV6m+fPjgClWhh9ugvTQT7pht
Dfz25jaEWhP/PVnZ4e8Z7IlJOKgq5WI2B6nnFTR08LN2Sqgg/vs4XUPGj2n8Y02/JoE9U2i+4MKZ
xb+sLu0t5fuMS24mM4NcDCw5o0zmUdC4D2o5KnesUBw8MHIkYnmJXO0OspTwMcDyo2mQWsb9u8IS
vY8wvcUGswCFRpP9UpFcmmmqHcENVmqCs/MEBEUDuVKlHzYiOyU/MH3mUcxS+Y8kp1n9dpJbJZ6K
4TuEzbOyJ6OGoNtvSZQwwAklmEkCqvUNRAfYpDBYUQrB0vEZLxs9lf1udUaEKl0RL4JBr3BMHZCH
dZHkDjmsASHqYjKgSYKUaakUWOSOHaVOfGa7gu0AxHFwNZ5dQONjn2vSy8BuoTC7PpsKV/m156Qw
XWor25NXccIvfFNL0M9tHzhVGaMKUNnc7bcg0ikKgUYo1n6OvwmMJB/DB7usbvnignSi+lTTPNrd
h0pqs04Av4faW4Ok/PI2PVePP8wNCchv2ClNa3WaQ4QMRATSpx6XwOOLJbAIcJwSry70EFD++pm6
uS9/EiJwFoGYcpv+Rc4mE9kmEiBrQzBEGgCkVjvdAY/B2ipqmUSDFvZYRXtLepH6tbyQR5/LWApu
xM1LkdD9AZ8tS090UjKD6ZEwghmrC2+gsmJ6adDPsttAk2P3fyAGfXWV2LP++bZ8iqNtyhEOp1bw
IbdZzQZh1bFx+tTkBGv3SYPnLBsc2fJVf2wgmPAxh8Pda7f8q90AKCj2nUSjtnGXZbDN8VTPd0Gv
pF7hgGpsQzmH7kg54MjL/dk1J/Va0JYumHcwyIYffMtWfTEu7Zm9h2iljbU2gwp8IU+d+vmNNZkI
SypRRHKnwexjASkzBEnX5d/LhiH4Gnun4ejl2spEjjgerQISTQl5OYtR6W8f7lv2c6jaOwO9qxnt
CKicRdnWqJkWsTSACb6+3jArlzRh9QvcCI4ibS7VBrsBpH1sjq1KwNbsf17jinnkpEQYSG+OMndy
2+85ISfN2n0ppn3nIsxuo+IO7dhlLcFDuYfD2aMSP/l4EY3syXiGWGABQZE4XnvWzXMivWCD1WSY
FsP0r4bkdgtF4rc9q61T0ssahBrR1KnEKBxkopP8obBxV/qb1HHfzLbFZpWCDrZWYneb1QswKCkO
jm4AJRGqKF45dG8Q1js9MfWh1o+j4jB3qYt5quwH1ll8/07nwGIAmhiUjYnzahAjb1glNCr8Uo0f
KCVRLjwVLVHSNdluQiXuV7W1mqyzy4vIsHeBJS6yHAu2ci/Pa0mpt5/DIMlhUhxZfUd1iF8Nvw5Z
9wQgDnHHTDIuBuJ3dE+VZK/OmB5rWbDLc4Xh4HxgsZr3E1upRjU0/S624z1AW3YglHaKs8noYgvN
H0TCDLNMUFlEZ5d5Ae9tkZqW8g3mncYGlIoHs16wi84DguHazYRGPmVAvupxgkj4IVySqeRv7/9P
xLkixMFRv0Kf1OeoO2GtK/v9FTtCQTKXQkJliUsbeLqBNC6NxU/UUaO3tKhdXDHQzBDKstZXzz7Y
JLAS3CsksWiH14p6ubjJkbcLUvL3HZRUxyJeypdmncvbyU1tXPXV0vceKll1rM8gz/fCag4Ar4T/
0aRHoDu239sXYUupjI57mmb7fx6LBbwMp22U1AxO76ir+WK2VwJywtAETWMndbBoI+iB1Qpt1/FV
rMIczbiU/T0LzFq6ntS32I5xgMKdiHKB+efmXSzwS8nzLN58tDTSoO9KeoRQFAmWGXRjK2dNUJhW
UVswlr4mAGeK+ZBYwtUkMvEbci5YVLfnPgyYh+bqAoInZvtXvbghESmNo0L+a3LpVbLoxl11vHWc
NAhjUS05abPWtfZIndTxhbmnMOlizUWxSpsBqIiJxp7DOTSNalw8Tl1Ka/qmDf2KNouQok7Jhba0
De/euwV9LKCbRp6NM0c2TE/dAaIlOOOcutqCL35XaXDRIQB2W4o2oZ8f/eH30ggjv9a1xqCmUdMx
vOm5riO8TyBLfqVWUwA+Cl9TLSCraynX+tC+VMxqVtvJrfmVImzzhHGCYEhYcLWHqd02M0pAp/+P
OzWkd/0oJ1vTAJUMZNK2Nvu+sB3UFCokaxqKqbfGhX6D9GefH78W3UBvMVYueD7z4vZOQGtvn5Vc
2k6R586pXc4viUEPOra9ozIuI6kkz2sMxRMEMAN8uk9wXVmqpsDEuXiK0Y+I2PQHkxWY0oFCdiPU
RmL7JJb+VYIszVz0ZUU9oq72ItyCo4cKvZcMSrGqnls4B1/dvqLWSCfnc+Pz2Q0+z7InBQmDb7Ub
yP5IcJMW57fUbz2n3uPscJRr/4OP9NxNP9Ytjgk2cqBae04xo7nIEmgccdYo2nd9xH9o3DwYKSGK
wovlufjcvEDt7vt0JQ/Hre3xWp9zrq5tJyuoMfdGWPlgcVTGA1TqMWcbV2/dPCKSt3b+aoxCS/zg
5AvOlBdM/1qEDj0iL+UzNgDczKPoiwYS8VKxHiieaK6eUi8qDN3cTEi3r8S4S6geQvBCQnInBF6G
KXoI0N9PmPslNznHxfu85buarRJWVZkhVwChEgpe39H5/nAuv52rV8XZ5PgbvxTXwCNT3usxNo9N
IW87CQ4RiFDGcqcaUKbpdQ3YBP4apW0/iPBMfuCxxhD8LY6mBnxegw7aDkkQ49rAMMdZXd+zqfe8
XklQJGFIS3xzKY+XYa3EXuWyyXELv93hP1qYH8zX9c6vGMnV+p7d1hAuN+nMxt/Z99VP2R2XbM4R
f3w/aQrzsM7fiEOWhWFb5XAz8t+ayR1lrDnc+PtyID22p5kw45HZ4+dn22JDJVrKRfrTWnQrTZ/f
ECU2fhcvhGA5+Jte0EflZf7xXHAR8/gBlMwERFQ5acj2FoLi94X8TeI7wliBgtefTr/RQG5653b0
6/6oYUmDYXcdNSk9Oz1XwwNPEUkN9EYtwiR8YeyIMElXTjN2j2zZj21A+PQxksLYrGbM/9y7cqJl
W0QmHvQYEiivg+vZLxyFYAS1B6XHkXSflSwd6OhXmlPVQd35uFW9/LO+p2kjMB+2i3vHdDC4p3lY
mCIApCNyxjbxqdLJXb3xb58yKNmXFsnhylSEAHS0d/EBr10KtpbfJCv7G4gLYlrotX728tg/pnOG
EZbXYmcoaw6EY0OkQFM3yqR3NFCMr7L+b+uxXmWR+v1l942zK2CLrL68PD1tJyymxh6LE7fUWDdA
Ov9LzjoFz6pEHWA2O/jlO4+nq20V8RmUL6CnVso/mdmjRBG3V7hnMTzEdIyK+xKqO2XsJeYyO1Sw
S1Knns+TtYqY4x7tuDm/qqiBk8TQUz52PvDBRa5p41rKvHse8Ut7+o9XJK5mwcOFijsOtdtBKqHr
dP/WnDbBvHwD8AOPoyo742FXMB/jkFBJoTtejK4HhmtfHr6hafwBTQCpQOZHdA/1OBKrfgGB8keo
CaXTpQl8TtRP8tsjbm1tKqVw0iHSfQxOn3IDQ0vN6objx6k/+n8EbWpuayx+SP6anKc3sf3gZNA6
9y44+kB/AvYgqQhOuel/k3GIjIvxVy3uAjtO2kGHf7mZw7fHopnJqgFAdE4V/x+R0u6d9qPCqtz8
ZHeDPNdw+Cyy2KQXftv/jIHZDS19MjGzQIPxo0oooZdZM7/C6Fl/ZFpJLlUlA8aPIjKWO1EkPEbN
ByJ50GI0/lmfTgHRY8dVGH2Oz3PHvc0IHDH9qQzyQLCIide9MEpzPFz66A6k5KD5u1NKNjhzFcTm
DxOnEV+LVw2xdQZaU5fwN0GXrlZFu06Ina54mi0VWaYn2LEZQnMiKmR+tNXhfYCb17ZO9zDUn58S
n9bHeqvgW093tueDHaQhRGzqCAOPhXUD9rjFz3/OSY0eEHlTPYjdMuKNWrMW+Ze/TL4W9ubRl+hu
rGj5cVUbJNafQhRKbuuCIGFremloqVboVnhyYj1yOJWXvmuyq+TRxBL+9aFNGmcDLcWTOu/YDDSE
nEtMLS4+T1hBDKlLWAiuqSKWQYF+MqfzqCfyVzeg1OSkiqfHzV/dscNV1ci527oXd460xh+4CQKf
nU9T/XM8Af/zIoPUllsZ/EppMUHq81C0YGBsoydTwKel6grwKD9ngyrhtO/TCfxnK/MBbJ5PS/WV
fa7ymTyKGRfVTZ6RqxPYehijPPAhDfRiuK2/cs/RHkeyPxluDGKLJ4Wk6IxW2bJv4gQK4iKbZqI2
gugAjofbPcaSWlfy84PnxRtgJc0hbgnZjWFY6FCFVR/sI1+o6a4YyQZ9mdz4o/MUhGkEnuEq5xJL
KB7YxFrWU7wnwU6y0RyjcIaJsKRQCF79JB5eEV5heIYo4C39RKZeVzxRnAHFLdSt0BGM5H0h8xLS
DuGVrcSPs7zgRO2xRgZVw2OsZsgkiK06IbnVn1KH5GPXYOvOlYTJ5ox39kTjcrs4aidmx1JC7gG+
N3awzYzQ9SAM2dYvfvTbcDxPrCXWQuB61qDWOtBtUgqL+zGKcmAeH3F9lVBsf/nVJjjNGsvdR6vq
iC4ekySs0JSy7FeBsal2JJ2I/BYqsMXYqEf9hFpIdFyL4fdOoxRdT9Fv+PkMfa/Dm5MgAODcSbmJ
kPvF+UWxBXZxbYm8SiQjFc47RLKda52o/y8A46+Mrb+usp0sy/5HD2zVi1JbXjKlqmcNrtfiuxao
clNsr2D3pJT33ioMfeo4aMigkKsH15BIyEC/Fpilp+GTeBS4tge2B2fhyLSg9MU21ezUjHzr0dpV
fjxqrmPM4exN5Ks1c78vv0v75Caf1O9U4f0OtKIcjRSBmiIiNiyU+NaXwTY5XyfSAnO7vYsoPJ8m
F5/40pkdcu4XLvFfQRfkOJ+WJK5tH+75ay8MiDegffbv2TFv9Qqw4/4/BA/3tnoOj+kEUIarDQnq
O34RMNLHcjM0hteBC4x4J8fqqFyqZYEVveSmDfgV0X65pRY8S4y7WGvbpHW08gsLt56zX+/ibOE9
X/LtZSxxg1isunS4gaGPKIocJhZ7OnfZYouQ4h/SNL6WVtSlVoqDKkICjc2seRCjRECNk3r/OwqE
xpNVz6q+n0yt6QIguLGZLXqgtEqqfGx6Gd5YEQzpUvu0J+yGnLgs7b0zggLVUHfZL0oBX94AsGWu
UCEBZraTr3aD0st3gRKKLaayb0e6FLethQ9YWu5whUn/VDJAg4Nvf8lKdxfZpScbv7/MfHT28Tnl
eOGmxGJN9WZT7lul8aKF2ST1YWZSdaa3fmZhj5WIJqH3IAC36K27QsWKhh+HqAZEcv3smMN+iTBM
MI8HAbW2nrH/M4eM07eWBbP4unXpWlBNfPAxbiVNfnqvqOsWI2BjMxBw9aCZS/L/b2/duuWVHsBZ
yMs+OUTekGsx4zxwj0ptjbyN4zuFqhjJIa+MGqvw220dP5yT+RFWzlBNyYp/Ulq8kQ6zgI3r+3XZ
nrHlQEXnzq1+IT35+F0Q5pfYUgORNQab7peticvv7mXTc0H+PCL2wTzEd1GHJ8bID6AxxfGZqlJO
WqPpeT+VxnVrP1vZNekXHr5yZQGFkA9eA3VBGaZAxP7d7MTIsaWAzinzeeWOMMFijJJl5m9fYhuo
gW5Svwa6loyIDrFpbl/WW0cTe2ckGH2j8d8eA5R2UpoCToBdQFOM+BskJlahDVR8bnhUjXJZQobK
Vwz887lcZ5sgbvec+UJTBwfBt5mVkk+mr6UeUsvpv+LZDFRlk0WSgbkcBXDUdZIPNZSrB7D3/5DP
Hh1Xz1+nQF0SB4Uvw8b/VnGk07XcPxPFDD0dqZjQ8GEbnJ/Mkp15PEC2aonhGLxMhZFnmn1rmCAY
QnYPDYZPLnNSIrXV/1vyQCQRXSvI0toi7y/SqOgkZY1xdpWvlRGGnf8eotuTfSJB6QJs8t56DvYI
WM3Qrk1wUcem0mqf/7Ky4v5dufYTZCuKrXdNkpUCvoS9Zkgj28ar5BLt99/3WnwEu9Ev79TXiboE
nDDh3PQ8HLn9d4l6noUkxqvhBf1s0VS4O14pIk51mId4toweoqlVLfYAq0NIb96Yi9n9yUJ9gLCW
ZaBeg2h4sejbs97+QUsKOTUBpBMLmrqLfyZ9/JJosQYAZJQI3/mZFWgpSYQmjtWDOgM/Y4kbtXD3
FU26Pu0FagtizJkEHpIR7U5aKX3kPHTGVOouJWGEI+eCaGG/XTc3ylbNrFRJ1OtkbB9mMeJm+Ug5
gZbExoJ/u2UeNc2MM5gVcr8ErYtkORCsAGSXAZqPvEH/NEPBtTjaO6KSQiWpKUH24O7CuEh+Mzai
Fp3KSTzMDmvcM4n6EoJf6yEIHTSOei63qMfsZ3dY3+ApPk8jm7C2laosNpJMiHyj26Ppm39xV4c4
mCbIiZKtGIO6yD3oO7+RyZF92aMaHyCDKmz/9BqJOXfEriOqCgg5MQlQupw/nbdYH2AGINmltFaV
MRkQrZkeJ9KjYx6C8S+w8m7+Piv4+OXXSkFZOr7PZTCYywyNnoOoTUBcOkXJpIjRSErHitcj+sPT
iBe8wxpPPanc3LLaJQ5gByXsf3ivWpsXzSc8wnF/OeqP0dwAW+IKuhOwb1wu7JM8iEATvyCehgBD
K3BFvVPCbUzfMP7x25KKKD+qE8ul0Kqy5GHGWSyQzZaxON0/mB6G51/0NbfJaDn4Okd2mxZ3W5fw
/hm5G2P+gdM/tT6VR9gv0U1ocCEc3/XgrGNEdEFp12IqqsSEag8dPAmRgzOtQQ9TYe6+ot/7ctUk
yVj/k1S/xg6VwftJCjf+rJ9e93LZXXHqMizTYwv5riFZMWmfh19dcoGMfe0RoupFE2kDa466e7zA
hhgT2TcsTVjUTLTz/5xmK5mFVKg4osUG6tf6Tb4eJSq4HKj3IGmNgkJedBn1yHCOW30Zh+h0TkJC
QEZlxZ6ASjALhboszODQVOI6EeN9GbK1/C0AQiAsqPQ2qurZhJm2KeU3nKBaiEr7DEw1kYcGcAYK
3S58dxNZ9nn8Qd6vqO5ugIKEoV4bS6QJBIs8Hy6nC2JgF78hLvuRWHWVU31GeoquSl1mAg9/fBY5
rNkkgYSyYo76aNQ/RxwIZ+VgH6WISLaqqODHTU4rwv0sduYKpDHu/5YwNUHDVlS7OF+dLNGzeacw
NWKoEaBj1vA5Ybf4tSg+T9b4ThEyA3afhBAIRD8Nw2XNyJ/0sgX+iMEMOZDszdam9yuh4QL4/iAO
K82B8KPZAsohhxUGCpY3bejH6lQGLnDwvwFS5l25ptC7HLCB3Oez6azyMh3wD9kUHmARS02gEprR
WAqjr9EfGblLd8tzjxGdpTsDAU8+X7r3AQndwExvR/LMPO34AtAhwJo/+kqRuPk9WSicfkmA81X4
RmSleA6SML4J7NSy5wUva+O0s3k7fd8nze8xJtALmekEvjT2XQ8TsRjZS/TsjpNpN2kF9SADSRoQ
lPCMFT3EYOnpmbffmADSsKVMuwnAXqC68wu4adJvmSJOhpeCZDXwzj/la6cHJpYdc8gDFxqYtxI9
k1St0QmSKwzP9In4hd0U1onfMFfJ67yxguwn3MR1SvYV48BUlPQ52bRMF0TpLZAZYbwWcu5WTxvm
L/4Z3VgJEJAXrcWMVcI57Xe3nDWwX4585VE102rX7IEOLwDImFQ+WUBnLGH2trvAFG1cDq36hbil
FLtBJpk/flrXHUf4+w8zzcLzq17P5BGr3oCcHpSfqVRla3kndljy7AdScjiOlr7qfe+0lt+8/V7G
mbfwCz9iVbyPIVtvQgL0hal38UfKDPVNqyKACirDZOkT439iw4Oxqf3LU1C/EAhIgau0Pcxu52VX
StxO/8QdxzwX67TqFZMOWDmKmdYV+46x+RVFll1Xm0kjcnn35WQWIJAzaj+Y+vQLVJ8TxD5tQaXA
N/EMNDQzKzMU986/AeJfG8shSbj6YoQTu637BHfVHAdp1Um/oEpPTb+K3HoTB2LT3nhR45mAgT2M
ixTeFRk8dvgh8/X2Uz6C6Fwra12pk3FkZBJQGARU9qKUCjO9iCz+wh1xgNnGAXcvpBIcHTzOKDJg
caSp8Uevr9l8BN+qGWP/RRXBf/ydPoxXAMgZ5/VD5U/8yygHWimjbEITGXAmrrO8kxzsKpC6co2o
AQaOZHPWHMXT9I+vDfpxKUIVP5s6dj9thBftErXc31DhPtUJUiU6lEvon4886xADqKAKoBugrrNM
Ny35sDyPzVUZfJzAiaHrZEjGuzI17aJdk05GyrypzNmk1K2PnkmGUzX9KmkSFtY/6ofSlwEiC3Dt
fi/yfX7U4zU4eQOWhSA1ZHwQRTgFEe4dVq4RDWzplF85TQH45imDgQ/no5NmyV1QQXTu4vvvEZy8
zoOvw+GEL18G5IiAv+hmXtczbpCPeVZJQjX3gCAw746BNjfmjFj07Cc7Fs2YtgkTgfHGh/wIpvDL
cJbsmal/Iwn8Rrd33R2aDO4IeErOd8/tyuAJmSBIwDx4vKvAPDMDmDOEJ11QC/Rrem9UeURYY+0w
b4ZNZmlFoDlkiuJAxGxAokI1UYjknP3YeJS0x0lREcYGfaP1uy5GICrYMOs+AflsOFLqSdrcgkY6
gho/86TgpKL1ioeabfOjp7v3dZ70ttiPVUQhFEx4stBEM+OT03M9fJibQWy7JiEi4pGONyndjYfG
3dfeM0EN6RdL0BvTnTj4PuZ+xYhcFUiwFdC1dmPMvvZYNWMFuKxFZj6Txa+iWvfiQ0gPLoaOOBm3
Repi5lpevPM5lpFpcRBGDtmS71woMh9RN77ZBSFPaQiwfCvPaALDKLp/2So8mkqRFfGrb2E9n+dM
w3kL+ZGycmR5Z1drILSItvNZczRCWjL2nQbQtprFap6W2gVNeFQP8jtNmLQ0L6M0QSIQ5hU1suMm
nBEKRp3zkYskA3z62SsKWMQ8GDS1osXoTfj0s30kMpEykSSyMYST2cvjQPFBPrxJIi5eyzDBvdMV
OfhpvQsLCjnqiLx8DpMoA4SinIXVFILY6f0lGDTtY8aEWM7uyzgJLBigY6HwFCiIjtQrc4aWXOh/
EznHxnjJke7pnsK/lEsW7PxUxN3EGbelZM23FS+bu+DxpBWWrcJzSX36vnWa48tNUT7NtmQaB4Jj
PIqwWv/Q+BK9GeFWb4Ubp/5eZjlQ8zXCf/D4jjN4OTZhYeUChPlHWsAEmoGN/QK3rFMO9f/H/yKH
/06+g5Uej74jdKqmEPm/kPogXVWsB9MqAxIC/P+ShwAZZ67ASqIHeJXCghYoa6q38ZQCMSbCLHM3
fDln9V79T63jGAtIf+EESYGuGt6h2YRWlMO8LWYAJbqD5WNLWEfV1BT3zvxSTw8ASm5V2OkVcKV1
Pi5XhWST6RiX+ehjQ7m0QrhKAuj9r83H8WmUbRmOxQEpBBg0tqUmZzJbmnADR8idYZuh3wL5KEn/
n0WrSS7TFKjf96aWyy7xfKTlIJ2pjF5cxrUEzZ9NQMfJ80iMZG04XC6JNbjjf2e5zYPMw0sCliWr
+wNaQLOCRM2qe7aEfkEgQULaBAGnNxbHiTJBRYR7xcnAk+Ewq63hjlQmHf7o3dkkYx9RyFIdMHZb
51yPix2VLyJqHg1P44OGzPHK8JqEnIUKgW+G362uphvsrYzFyT/X2uKXrns5/tTBNQzxrF9bsngw
J6tRKDHVhAM2oKBLWX/Guyrp66kaYzwSG4k7uR7j2xwvEC8OHk/RqCE9BPeK9YHGW2hKNjOwfI6q
RhiRHblxO6V9LpWHUiQlT0N/300SyNERVdDSteTtNsPw0zDNL6jlfQ/opi/Qj5jMOsghwvRaIM6E
TJYzD90ogW76zQSXepEQ1HntvSKJcuB+hvH84GbmxvhrjNyAZ+1AwkQiV2PZ2Jl8Ec6TMtBJieVP
KAft0tHmujgz9XdN3hkdKj2zDP4GFf2Nzw3NMimuL1eeiyprsZSSPeqBC5cyw50VLJGBmv+7j1hB
ZBLorNr1NN17bl3BFgSbOn8ISiQu7HPQU2EdNjgaGaTNrKQdv83xWeIeo0GDq2/TPCaJ4wZpSH9Y
P35JwF/XIHgio7HG+xq63eIiisflmg1OIn2WZ3b+1rfw4WQPgBup4EYuB6TGXtR05ZRC5axUwtwW
jcS72Sm9BIuDfOa2lO4RL7XRB6suzYTev/P8ZA3kFrRpLUMt7Zs7ukz/X1MtRAUqMdMXi8h17hnU
k/UmiAqKQ9/FidPfcIlbmckb1YXRVibNPqv9GIVAL0ORV/8zHDDc/bU9d0FmAX6Zfeoc1H5fRcrn
2/wv2Asw+SYkrCaVQdx3x3/KxK963AoJMnSEbCjqj7JcSRJVEqiKbJWXkgXUR2DfkLSwoVEbK8RW
qq8FM3ugh1yA3p6GlPag24ai7hhlbQxEMVzgPkQ+gjB6BetxdzPWnISgzOvsMyZtWrjqDYFq+AtB
MJOTbMI2NWT7Ob7yTBg3pam+zKuksZhmdlUEm3T+F5lL/lLbDlj6060mC8hwYTBMnq5+Jh4Pa54v
WVr0ywqUhfRcYitAskDiWroHC4jLrOBCQQH9S2FnhlHfn3zORTNrhAA6Q+QVizMn783REMLtEvaN
+A8Jhf/ftUrk3qE6fIoNbk8NEfjlIz9/O9dn7sgg9sdDFTiDs6TzbovSidIxl2Od85tk51l3Z5v6
fkl3FKQuhipDsQqAggvk/TJ9WVmN5yEVbEb3CPCop+xKO3wW8BX7WOkTiHK+Z3v1N7dkE0BHZ59n
ZP4+7UzJFtIDEpgEUh1Jyc3k2QP1uDBRaroGjWUEEAxL39jHWUR23hAcHFlH9Ogn8uk8Dp62lOl4
fadxuSaQ8Ry5+ZdzknnJHqBRlf2xPgfBs9gPhWVz7w/ROv3tPYPvyMBG+UVMB9cjxeMNyZLMkMrN
Lw9kAQjLGAtBctRuMs2ZChPGKylz8yaPOx31UqKaIpBtFqFT7P8HrV8Pbpby4aiYeTp+awnVFlCE
djG2IP0UvH6pctUcfWSDT/sETxziKRGbAOrKn6JNISg43LZv+B4Oj3onG/EE7gN57PkrrB0RdXBR
MwRs7fxwOft8Cygy53mpGpBWBdvkIGvL8SDDNwY3htO7m6VLZQp1IbttGTzL/0SCG5QTbaijaqpi
5gjnw1ek35nnnCwvB0l2SGGd0YNpAlq/LQqTB/vCLUcKEUEShquYEUZL6BLG57I72uiZwpk9Rm/7
/YvvKwxQxWlzV26gDPD2oSFvTA3NhoPHob5XgqT/cKJtURk9HyljE7x5JM/EMBuPGuofSSYAoIJ/
7tT5HjeLHz37vR5yr3l5HfXnv6FbiSaSyIo9whLcL9Ote07yrIZoxoDl3pMLkC2fkgBbCf54x3ou
b3KngMQD9C7vg3yfx1ysFqC6zOjHAnKlBPvxmYvhOOom5BPgsIfWlS4ZOgOf/fvhSVsT13CyhoRs
Px1GmcSUH3WKCrd+aviAuaUdP6ntgXzOwuv3ScoGa0eev//kwe9S516H/70XIaSFwHVNnitAQPyD
Nd0UJ9N20taElBjshJpbuCJ4jA1uEQdrxlbeR2ahakaXXc+RcsNljfnSo0d6ZQ/Zuh7knNzgW+QS
23CF8fIqxrtcjmocX7LMaxY5BhRr920/bNFPDQjRZeTMFDsbt9L+J0h0bql+/eQuc4WJ4OQicvi4
8QK54Cxt+Ms1LoeAOs55HZUjMw2iKtw+zs4LjopZCfhyp3F8lua4p6TTfYKmzhCeTnwMVwpqk9Jg
kwkzl0LEsH6XJmt+U6Z8aQ/EmJkkM3PDvyEyn+gla9E+tkdjtch5BhJehIbmm2JRMM+6aOrPGLj5
XuqPlbTJZbiQgAUg9jWEJzwCEE27dsqGAmmQUIDFFLrf/XROkc1FjWuVVszdzdf930XTBl9fvvTB
0f/g35i5/piehP1vKGylcUv7T4yXT25/Umz8p/WsyEfoJ9VU7mbp78AUUL3V/1F/SQ7pIEpRoT7w
RBp6ZRFrJh+cT5pagEHFVyf7v6KuhKrziHAYDfhSpsqNZd0xhd47yFv77ol1ec7w1z+SNnLLasy5
OlwDFAGDlYi9pwHOjeEZlAM11/DQlkGJDg6wLlYXj7zptwjztCJ3DOmHG8CMh3N3n0vKCYzzlEEA
cN30aLkC7BY7cLYHNNesKRbEOJhaOO4fSMeKTKKyQ/A0zJbARoiQ2dVJkLZYgwMAWysy/RsuLO6S
ZFAuFgyx9USSOmFRBw7/PexVKG8SKlB386fAJ073v1HCgook6AdKcKMFwZgV0a31CegzfBkFMa1g
AapHoBuCaiU5Vhw2Loz9TozXA2VL07DNtrtyAMhguijibf9cyw5GuL23U6+9yYj72n5+p7SNqmnK
qW0OcLpaiNBO5X5vBH82xzWGAzMYCChtidq6I8KsjKsmUSM/Jpw3JpEgXExCwiHxwWwFWp6zaxmo
vBkdLsm3Ru6YhX6ZF8/OErTb+Gzpf6GhsZFGcTwRLC1s1wRwe0qd0HiWdsxp5vxVY4IOmAFfII/L
7W5smNE5CexF1c0CCJZ+mRots2B866LidQ+KNWnuA5yLy6hvOxS9zM28ZurvllJ5DYnJ9X9QwXi5
cg+uaYYDbjeW9BpHeVmAIFLrgS4y0I1WlCtQZKm3ErvGVexPd0gqkMyQCJaiqldLlRMypOcUpG5r
jtkpxhifPSVcFl6e9YP9ZXnfN6zOAK8F3F/NdEZYnxz5WMIB507AjrvpM7Bu8JzRDHsR+c2ZWbMQ
YJzQkKp5sBLqkEtbiW4CXig+V/k3mrZbsPG/iKpX34Rb23Fy8W4FYhH/DLzTfg+HEOtpjeB9wLbu
iQwe5xrzKLUG1zQg0K9nm6HkhfnWUjtFN/9YKiLu2Ze3MD5h306DBCHgU5jC9PzKgN2tQeKhO50a
j0E79Klt7M9J+CZf/cCeAeFLfAuBYFp1QQ+J5Fac43gDaDriDAWl/1AtJhnCKfs1UjcOQaIp8GxZ
a5OasXr7iJgSm401iIXopOujxsdKS3dVPB4kucQFRTzbtUGremuhLAzQHLqsDhQC4cyoeVqR3Xcn
+y+tjmBArrlEHU7uA5GPa/ePBv88wzyXbsZhRtWX5SXHVnoEChvWxsHunLPSgYuGYKrtApXorDQ4
py3j4kW7crsuCQ4MGOdg5WGRw3BYy4qUvt/qqpXpZ6fptT9foQf/qU6MrxffxeIS8h0CHsmPQlcx
721spfm2H5Rlsoh25u+KsrXhwKkDCupA1Nivzr8iyEoofna6H7SnuXPAxETbaxCrOhZBI8yBc798
BbVl7VUsaKdXeklXczTZLX1VSCkPPWVXEfSTRcpsINAGwsn0dj2pLygYlB/adxhhphHVaTx+H/Oc
RHMTHSYwsabHg9pUL+GoLFNI53ujOogx5wi3WuLFfU665U/g9zPCfNnXlOhB6kQU6k8HLKANYU23
xtqHDkCTuYgtr2aDtPoJE1baxgFUpJOhd1KNGWjBK4h/cDCM+HilrXzDgvOhPu1FcmdvLlZnA4js
Tjx06KPDvRe77N064lXGGAWHhK4C2wLNh2vJdNtJlK7FrHf5e1ifTzdCdIYD1d8JKLYMLbwCKfoL
ToDCd8yGOwamU1OlGOgSNn04qSmyeuvQRYObr1yWL5SdN1XgYSp1ZUJ17+orAHmC9JWJ/4jFeGX2
7xNcapBvdTTnldLteg91EHujjcKznqyCZzimRAaxJnwOOY+S+xhtte9AXkHPMeY8MMTxz7iNxHmR
BAh5WyW08BMjDhNgFY2cYfVA/7MugqlmjfQMGHwAbTPJF81nvn6cjP+lHQ6CYv29fbJgDWDW2DPp
aAMDNudHOt1dz0LOqmC/oPc74ee2dsHTVaF5TUDlGjchMBPUaUICqMQGe2Dht+sM/ubM/4YU1Ig6
eoh66rWlqXku0Y/jLa03Fk9lQIhYHizNoTDuHTMczEfKawt3VH6OQWv0oa6HnHFPMR556XZFS2Ff
qkxmKI6MtISBk0HtiJAilOuoTqbqcpUDwoTRVrt0+w+gUQUlHW9cg5BSS8aHznjQDDzwH+nXPH4g
7ASKlecWYG2USbu/25OMtStnS3cbGPc8ZV0b9un4DoykR/WhmADj7RTETmIuVt1rMK4+gfnQqZtw
/xcecoU/5K+xD6xOidoV0pAy6nmt3RrUmOZw3qVW+mIGZBq/x4uF464r7c1LuyDeMrlg/atbgKA7
710yut9o+Yfi6aF4ohi047FbCMiOTs8QqACQuJT/NWh2U5nVNVXX4v35ZHAY5CcPXUcSen9uuV68
qM3ZOmr8slgm2LTj5PM3Zc8mVl9oPUtgj6h1TP1DsJ0oDgAq9jv2T7/cMiFhl/6Z2QygMftRw3Re
VObYr2pf3qJ/MNaj4ErUznT3eR+cIk+RFxKmCm4kvKsUNigmQWhrRrxyP/6HUyLvfSLNkjyUUiCD
M2h8zRz2u5uUSTKCmIZSZhV6+l8u3O/RXr2RDVvs5YL75hrudRjV00sW2ca00NH3T1dpWnJ1RBHK
ysw/m20U0RP2hGdqZSY1Rb7Cmev9XFCUWT5/ci7CrWX7UPTTkiDxZmt/rut5pd8jIGKIjHoUDo6e
j/ycCQDvJ7KzcKhP1ObzeInAId9hj91MgqcILCWD8lHHXHtDb2IwjVepex+nfilwAnoXS2BfjX9N
iwY7Z4wTsRyVfGnKUmwbcMugiMYM+KXouptMKLdHOT0+5HlMjkIMgIIN9oBone7b+fAYYU55nD9b
7JElNhveVhPEXYHtUSk56f41LhLG3i9aj+iGAYpMJbktw5O5ziBjYAxVefmohqmETqwnkGCUSnU9
rJc+gZmc1D4NC0spakJxWPrbswx/5qCaPmzPvBuELuQdKiLblcncLsGLhqnZz9IRR8DdkLcUAcoR
EY1eWEG8Eww6bD+DZdOyb8jDK05geINlKVD7Z4tG5/mW8iYp3sa1LwLQbPBChoLWHuNvxN1yS+1n
Fv3i7KLkUQrz4Dn8unKJy59iqKUr+wN6kBzUHkNX7vTh/yM9Ke2eY9GM5ViIBadmUiwz1v5y3fSr
5fjadfX5jbVaJX5L6zGGeFIwsJTt7AXp7qGrfimdoZp3KskVr6QZ7tpJZEAD4WP8ARhB6Rl7swe8
oy9mSBokOO8nPgqzwEOYwfGTVUNIHsxSVB1AD/e44EH2RNTCYNuPdNiyx92vcappYTMi8fkziHLw
NGpL84hUnFNBCoHZCk5/w1eqfSXsgS/Xe2biUih9xyO3uXzp/ON5pwyZ1WuoVWNzk63+u8uUcQoI
hT2PFDDMM86B6UMgcNpl+cUkuDHOSlhIAY1wh6Q6c3kHh3nVeow5sCv2060M8TFz1tVYJnYb60/V
WRHDj2PlUUChSh++XNam80Z+Et9SaULm+xsW5z0vKA0CB/sex2U1DSIiAttnb9KOy4OHmY/snL2/
9DMXuumR2DZ382MF+M2iO7bShktIPqZHmM5xWxKHB65nwhZ8alsAIzV+tjUk2gnRxpiCHRmosFQq
SxD/yjc+f/3KsshtbYavfpjN8wpSwyElFk6atKU48x7LR2CT0fFrLqfHhJACn87wqBx7/1sPZNrw
DeNHumqOIJ7sn4F6cYY11B2eO0SWnXLT6FkbyVzafZgiBzOBiSxnDBx+PQP7dJtJhStsd7NgtUpj
kzCflIZ0cBS2mG9Jbqzosr3HB+3Uu0dBJ2x3kNmJoImki+npLilPg3LDale9vBtsFindpg/RHuPJ
3IiC+0Fe4wHGqk3ewGxtdJYdgcP5gq7weggbUTlhhnYVixZy+TSr96JAb+d3QU9NimyCGBB9O2TM
vuMtDvOYWk519JQboChgiakT2vZt8ZFvmlUg1Mb9LfOEGFzb0d6Wc9SkFVMrN8Y80FrSDpuKXqKK
70sZT1+MaDa4XH8Z1fL7SDvZDb8LZJq4/kBGeJLdL0HlbXczTFxrLQ/6DZMU4FdJv7qMilUILNlQ
6qHKdAizN4u+Xhtz+6NzObqlmld5Hn8K0uz9e/IeM0Iy4Ewg10nFXEp0c4yryDtcMgD/rHOEwH7V
o72qMya4XquvUHn+3vgYga8A5yuaMlycM342ANtPInpc+BVJDhi9mySvLX2wLPWhoZs48B9nlZZu
Bgv6a5od6KLin/DlZavKrs+mciFxPT4QBCSzh1gjPCScFAP450jCxCjyBuOE+pPCdnBSPASxzye8
JaoEDt7XXnm+dQ9wZHWtLzrIA3wBwpWpSsGl+oh0W0bnYGK01RPhwiWxXeOTLmcHvcSxzU/pkbnN
VS2pjydXSig4mNt9COO+EJ4b7+qsGJgKGnNKQ9ToNcGO25xP83Gnp2O7tchlUUTrhtY9Wf+lRU4R
pXlFXQ1qu8+L1jzTeW1F057ONrE6v8SgF19Ix6stGbg1qACKFEwYYttiP8fN8/qeVTO6L+GOlozq
lP/MdP6qfYccJvHNMDyjbNPMChCJ4YmRpabal80i8bNp4kbyNzXZuknZoiF39cTKzXOtFefF43lL
N7ggREemBdjVF5XKA6+kfvOa/2VC27731b9YusjFOh5WWDessO/A7Q5bzohx+IJmTilbzrniFQC4
fej1Yt7x3s9MKW8c2Yx5YE0QZnH50C4XobUESmVdJgXcjLSkw6gTdRq7jPvkqIiTB1CudSlgVtS9
tJCV45fnCttLOwCrfw0Ld3D7FF82QdTrgjVMjGUr9s9ka2Wv0R7ArS4MkqbEUv3+FSf330wqWt59
f2xv2JZ92Vo+U/58Kqq9a41nEjv3Wk4po3m/1rXmEhIRnvxSMBNz+hu/QyiyDRiUk7Hec1RMLrV9
1r/1DP9mkgWMpE7ABmkHG6SI/rFAKn2tHNp28JvxwXqT082+NA+Cawxnc6zEDF8iMzmYkrAIRT7y
nc1TVSyRkAyhBrFTcebXoTXtvZ8LSGdLCmxNg2Xu1ceQTi+fMgwk15fbZx2uRxteKlHkhTUZttFY
c+6fTTvSSBbvu+MbqLQR7qkzfetNcE9d/awBtcRPrsf3yR6BfQloM7fFOuCAwourAqKz+c3PNqcm
CXLH8gyUSfKMKXnGn81P3eytcAdyyKpW+YYncIpM0TkQQWQJsUcOD4biXP/RgPKMqD1d0O937iuo
rhSw2IBBi1IOJ73FnukBV6IppqY44fZ6HVicudrkx0KkyLPijndZ5poy6qNGqDOoTZFtIx58GQ40
bNNvu8EV01LliLOPhBuwcUoBvvE0Kfpk9tfaAw0QN/z3/KDmZGTiyfoBL/Ymm6CTeRXhwGSdk99P
Tmyy6A/3YKqeutsVebwiRZoVKW6+b42idkaUUxMN3a3l5sxj46b6EzznNL0eEH/MoBWXEnaGmw9w
oHmT+i69gkSU9p2tGUILSaAUO8iZrjSYqEWREGg3VtZhBJbhHEtnwGRiQuE3wsrKE/fq/q1X5uiA
eyJB21bxbL1dDRu0oB0JCwc7Akvkxrl40w+vK9wRpeMBSfdGa5LzYf6iyaCA5EEZr/DN4zB8x1WO
ZDEbGN2euM+aGK/38lrUSXlyvXmEHQ0mb9aRs9KosJXfrhi/feevMkOEr2CG8zOF+6+I9wEWBAb2
7QSXlFSf8zJiFhEgL4ARUbYxZmcznx1+Kz/aR+8jVyGcG6rdyMzyOS/JZREOxHp4bxtuH9RRdvGe
Rl3LEo2aZXMlJpqEUgzAYUDn7yM/QjTZxAP50jlAWRXkPyymGfO23eSBg1PkNFMZpnwUVEJ8NZ10
HyNdpFxySVdU7Ht3Kb+fUHCZ3LCq2OVviG8lxRQ97xim5BDZa72GbxTE9cOKNNwdD/J1z0yP4PZS
MAuYm/cdQBrbmD8vN4fr/LKPbS6DjPas4DdtKkxnZFr4AXOtTxn9EoIfUNve4eLI6Qr2ecsUqKLV
BA2DOBtaN2qo1BO7v5e4UGe5KcpogO6zGMBO81mv/nR+/DjpzKw5BMFxeKypBxZ4TCVFc8uEfRHw
+0BPHDlt1IiuKy8spXfqriE0eeitrOYJk0zDh9w9D34VmEntBTHS98sftd3ClNBrFZFiHGBmHkg8
rdxYxMU1vgNE3Gn/OB3Z8sui+tsXF7YeHrjou2u0E37F4FLrE/EUwzsjplF7M9MqNJeFaiYZO1mV
23/6gDCSpTz1y9Z8shZiVRnv9vEZB1CZ2rBmXKIIr8KG8KP31Nj1M2h2H0rLVP2bEqlxNlzcZaNO
jD7RI6EfSawU+mpPNAwm9NhkRup0Hi/v3ClRrR/JG2QbyreUeN6DHbBSoDKWCQyv21QnwJVCdYHv
SS0yNWeQSHOT2KwQsotywnUibfnmUbijJSMzfrrEOTTIm+96SH3B30cUbkcMZYSwcA8l+/lOb1e1
MxjIp/zT3ctYFRw8bg/t21yG6nkyfwB92msAEh7MOB/Wn/Zg6+vMAcXQd9NLjFFOltX4a58v7RUw
TbFdy3q1KHFcETvNNDKhZCLy06w3ebpzbzLHfHDrOrvwQaUjYLMgnqKNClAztoUvn1FMQP/Dfr/6
EutIcGpn14rZE5gy22rysruHLgNjQa+YsJIQ8Dr8m1HcB6P5ndd8alyCJAxPbnPIgXoWeZ+xuG/d
SxZnaCLvPsazP2OR7zBdHHfl4yPFbLDSzkgW0g/+sxUXCpGZeqmdPpUrdL7Rp/BZmhjt27F0xA9D
eAFgk50RF1RBptP11/IScXv1cjXmXH67wquZskI3TiqEtaLof+PDrKsETlPF7JDyNAgTPaC4x8Pl
ivRO7Gcdf0AF+Myw4+xEr4gwXbCt2Ajud6ZZvNUliC49/PV82xVgfgjM4KZCfxONgNmSrGlMTobI
N4vjzNzwRNhKqrZHqCi7yZNNwEDpwvOjL6z5QvLk35SI84//tjzfwoEB1ZVUFZwWzC3WV2Rq1iCI
xN5Dxv+8hDDH0xuZ9X1uH/1SYO7oDmiUyE8YjHKgnzp9Wu46em2uprwJ2u3qePcSqcw3PfhwLgWJ
QumBnZL3sBu+H1ZMTzGdBMzOQ8qlMxqI/fTKfbjnPEP24mNSBnK8LYB7Yl+NcXmsTdyeO6Ic5411
mr4E/i5o6ScYipF9ayXCylgUEk+1LIw4pPeeS8q9fnv7IPLYt8iOGTDrqskHue6eeOw5x8COON30
6i7Ry4mctD3ppGc9vaCNdrlrR6AAedi4/TQRAXywYmek3YnWTc6cWkzGx9Duxpm7H2q9Cssn4GR/
HYRKJFZIcJqHmI821kFT/nPOpaS25eAsd7hAZZmNvbIU2hNqol3iacdpJZZinzlFrNELdLQPjeBc
K8hT7DBuC0oa3SW+TEmii7WyjV8nY6WaYaW7pg5il4HEo67XjPGlyW/dUCuLVloOdoM/5bbtEVfb
kOZdmKFGy0hXWf63ltoqDANrZAafQ3alrNvWV94X2UMKIpbaISyZHsS5C01SYXzTjEH17HfYlvHh
SN1K5/ZZ9FNFYbXsy+jZNp+DS/yT3Lz0vHhgQZRrTrxhPx+MiOJlE6tb6YY5XixLSFangG5/lxi8
cV7Xd66cUwreTfn4wU3koSA4usbbg0XeMNAu8e63dsI0NnMoJk6Fzf2TqMWBu3em2cTqH7tNmsKe
KV1Hjj5toWd2ioQYTaoPXNZXHXonOokfK7w6o/OHkdNHXh4LpDR6t2IJ4m89sOV/7PyEpPS/uzuh
IUE4ksomRFEg2w3pQyc4gpZdatK93JKSOCUcjdKWkbWhJSmw5ItGzwMlGA31m73OO4UELJ77TYjV
MY1OiDDGz37vW1d9Ax56MsYwaFZARY4wOfPGNfiyYoz/5tAQZZfjvbK3QWlduFzUD1QPC3BTv/5o
+zg+jtNW+U3kcvwXjuizDiKNUgZ31S10nxHX0Lj2CIniI7vUoTvUL2PmciyVdquLyp6fZgfCc7c4
zGA7qFqUVipUCbjZLxS1EttD9f5eoRC8q4KwVTM63km6bEMhy5/FPH2HK139GgANQMrPKM53D/H4
P9YaDTkMoBzNRVP1A2m+PJaLYHl0HcRmxOrMhAzhCPOR0eexclDfIHN95gae53AdO6n98f/PPsxA
pH1MmxdHfIWSUEbLVWn1xkSjLmKNAi7pxVn4mPgcnZClb50TZpcI4BxLxT3VsvaPT6TsktxV11zf
Kaf4cLzZzx/LJVVGZ8ZW3I4A5m8fBzTIlbWKWKgvPNu47EIdFtL91F/RvCI5fzjEivE53wuYlKQn
kxLqU2hWivCOC2oAw6IL+XxMsuwWhoF3zecLs9waq6c3OBgXGVhYxQwFITtGnUiBdYxd3SdkmBu8
PPlo/kBTPIPyWUZesrs5ZsiOCyIV9RcXAw5FTrHAQtFsCbcNrIgtBmVySbgemvv9PGbYXh0X+Ezg
9OHOhQzt5zQ+beLhkuaGe5Sg+KGb1n3JP35pvLY0eF3t5k0uXGx408DH8sbQW0GYmrkUHXFkwBdH
0gXr4GtBhVrkF56ZL7rNyNNCxszWlrykjTRzF5lSBYuQNniJ+24b1aC7hXDp+4HaFIBfPdIM08Oi
3JG+FYXY4PlFw8n8P9mRtlI97XZAISLu8CDzGua9UrjGGWONC1h7WqxgCTEYHY67sT+zYlH6ybiA
ndqcDyEO/YB+18vxaotuT6CHyZvZPN26B912V159m5IZqz4IVgFexm75iaKpdrkDM1A+TT3Aq68R
B6D1QpKn1Lxzt+VCEUmH8GwmTFRjFubQtsFhUIBpkukiLNmsrdfUunBUoNPlWAm2q90CDIhjAY9M
Ty5snean4TcpASV57b/WzPqTQWMV2zhny5e89pfFsZZfCWBJGwsK3N7gc92CkvVjiErW5NST98DW
MxeEd/E8u5mnu2Eglh9uoFCUhvWBDFzCGnkHtgEqD0BbxNpdDyVgguAybAfkB3VB5DRkwIbZLrrJ
eaWsI3aMsBrYdpKXsjwg4PPxGVxSyQEckkOl7691zz4Yul/PxvFMe/btbaUAmstOgZlRLbanbBFI
uAGV9ZKVCKGt5xyZe/FUFyxSoXxAw9fO+fbVXXqB7F9PHk+AXwI9YBLwVwGVtie4kXVvbCSjobAq
1ObHuzxx5FcTaQ8Sz7cA09CnSFtOJbjql1h0ufTROLp0j+QmOHXTmPYYknBPzqRY2cCnMvw70hWc
j3TkftANgyy2yox+pN8woWEqqgUFJqRGoFFxHn4XYn6R/p4/dQIeZzHYxeH3Aq4fefJsPO4zwMnp
YHTghAZzVF59+Z+9ec5gdllQm0Gmuo4bd6xPpJK1iDUmfTMQpfg6cEEs+u4a/2gAsxHlOVzOQwwm
ZCNVYLusn0cLIQVg6AbQ7S7yHf4AGA3ijNyrWDvjsMrEfV7NdQw7knVpK3/fEZcbjx+LQGXGh6RT
7o26oDNV35eW75cEQQW/+9LsfC0o/oIM4klRcrP1oC7UL/NpWmXSETpf+TGDMRqWfczzRUwg9rV9
fl4ofRO5piNPNWnRmlWTFwhnjV1s0fvrfxK4afHf+GBd7nW1ZJxk7rwsRWvgfq3xdcBuYsH01owF
rbnuWbBAklFAiG69aHAfMep11W880A27gDaYxgHgPWKdjmE7FD8m4UXzzYIIx85PgJjIDw87Is57
NPC2qbFrf06JLWK47SfR/29GUMes1017rzoQqyJLKz5AETT8Hsy+RfADxt6eUK628YYAjnnr9Pic
belM3AkRfruOaJvDtuohw5z8miQ6UlH3DlohhLvEYmXwWMwvOqI/uYj6fSGA4sSKZuGDhQxfBijK
JFR1x08A0RzxM9X0PSXsNQaMk8PQ813TFkl6pg5U0BPBWsUDTXrHBREvkfqiR6NCnGV5uAoDKu+O
2ZBsko8n8GSEh28SOrVj6+i7jkq40OHGy4VYVMq4fo5kZlKtFRbBF2ADQ9ZN9/r/4rRGyNlgvKCG
89frosPwtcRCiRU6fg9QTHH7SyLRwSdkTUx18rA2vqeZY3ApwyvTRGRbOI5vMEzFgKCMhxKR6p3Q
4UuhuIWh5Ee7kOniaH+kYPYD9OVwT3LpbnUlOqd9dDpxo/rtnYeSTEYXbyneOvAEBzwA3W+DyHQL
HUORmekL3t6It1uaXuu3Bm204qUeOL2vD2vaoUA1HdZgrAAtuNxc3oNilJE4E9DnnNkcKKblua3P
+BaQ6GqowP8yhSNEzcmBQ7Wd6vKa1Yu5nuA8Tivqjfw6tigpMh7OBaBJEtSjQA/ts3666rINZFpK
rBQJo9mHyBTHp1z4LX+Q4sZxjzUutd5/3Mu0cbLRLBNq/3NStAXzor+oyCQ6t2X9R+0dKLTzFeED
gjcOuiY7yzpyDBrYc52FmkhCQWjiHxFi1rrp1WFhV75uuPQ/gb8PSdCnMtClC1tW8uSpR/VmwQPP
1AgmiVBJ7BYOD8xZxhyl23ggn1PBLq2oLjJC9sfuwaKV2YbIfkPrI2Kkt3Wf820XK5A8WlkbEpOF
KGatsBL6Ob4Flxmx1sfAkqdyz3i21X9y+nqfI5Vc6XxRrDoxXdoC2ixdXhjZ5Yo9TopuK+i7j4CH
boPuAKwhqnDhc8ou63dkJdjoVmhiKhFCgQptekxfjTfJysznhezCv8LezW9nFiXf94bZ/fAvcljG
MoSpKiWaYyzsx9ieL3YTIdwE1PqTFKml/gYsV5LnYvMC44Zda875E95BMd/AkEcmzzVpT4z/E4+I
l5N32L9w2pHKag4HwLLBq2OPsgSNydc/KTrgy7ujTzzwx1t80PVsoASQeydVnxAo5wB8Gn2ef9+A
nJTZ/G8wuk8jWy4oVckDmLCHdD8f9ErX4K1y9oY+GNaWIzV9Zt0DFhWtX7nRFjEzJPMKxa4XhuLs
EmTYMeZ5M90eZS5X+lv9KD04+LLjPzNjkPU9CQ3+RKeDXISkgBVWc2RLFlTHpBw/sGA5DZxlaxVT
xy9sjpfHhQH2scRAOc98HJSZ94uMHsNIlE5A0OarXshQkl0SltOqKtlCeH17YynFyGrxnpGRZyZn
NPrN10R8heNpIBoix2pn+5CWAv2YjDxnf/6GIk+S+aQhOM4PXLCzpWcKEB4wCQR6KE38Whj/Xiye
kOuFRPDsLQ2bhy+IJolyEn9P+y9QU59olHu3QXOdnevIhNtGO8sAZPwVJgtru/9DvrMljkpOv1ps
XDTBQa5eWTcjGXzYlM/ahhAVuLQ0QoJRt2I9j4mVz1qH0Jl8YsrytnFfHcSdK5tKqFzcXwVNQNpq
cE0FpfbwNYL+pVJAKrLVyK0tFq8609gspAF5oJ66M/KoA0bkv3AiRCnBdq2E67+MF6PK/melY/3h
icMSgpC/QpsFa40ZywkbwVaw5JkHCpotrwmOjlEAkRMuUG4MXLGuUr8pR/omB8A2/x4mSumNtRPb
/AwIznoRB1cgN0LTh8T8ZDgyOWXrAJh3KBR2JDHSVqsMi1IHaVBWdHI+vgQqWD03FeQ823HdaIeP
/4k9xKWQbf7oKQjZVV5kzzvWKx0H9cOMD7ZHFO+fNONbu317MvUW3rW+RxY6zNobB5XtfVjmqdhz
cAgerz3DzLtQo8L+jGIFQzE33tVEnfKPk/gfeZI0lkpjZ2nm5vNFu+bYfliaOqNsjP/wKqI3/x3O
1FTJXQz8FU7MhkG3Hbvp179cKw9Ptvr2UK3UAuizlmmnB42LwnN6tZPl+LFPOGJsRIbvmNFxhBGO
AzUGDgbQqvXMCH2kkMyBELVNidBWBZVS+JmAKZMuPpw4drkuvehnxnWsNlQ0FiaoNs1RcvmkUYA6
6euQYOn+pVQBTFcEbyCSwFBPcibZ/wuT49ZaX7j/SMEqFzdKXAC3HuuEAM7awPSuD7LhaTUDrh1Y
ko8v7MjmLzfCT0mdEsylmBxVeH3fAd0pqlgRLGm58ksZTBnthJRzGlwNpAKFsKUb0DqkPrmPsxXS
bPne4Qg28nksyrwnIbg3d7LwbHaJ4BGUzUrlh7sXTn1JscuY2hXAWpZm/T7n2j0hhA8RlCYNHVPq
xIZlh7itwLAzvS245Zv5AhwTQvUVHkjknOcy6TEG3uVXb9QqnCuQszoeJO/ZhD4fPbC7aF9frdt4
zj4faKLqydi7gfubld1+M5hdmk4e5FgcfE1Pppp0rF4UE6ToE2TNujUFFpCa4H+9GdhZupT+XBKV
D45kkeBf32oGSWtu7dOgxwzYKLe+m9Sq1iWQgWwQBbCrf6KNXAa2VsNd5WIpr1/kdwf7DFmNvekx
1IJkwQxS1IsSNndZIaJswtErEbq6AONsdY0ZaDUhzDVSxxUYI3mMt6mh9Eemqh95s5lV2T0JUtiN
abOj65KYWD2amEACh+ZtOfOrW4cwVXwjvjoPNUfNPrmzZ7JyFv0rcSGiBkMMpvxSN/1tNteTXdiS
vJCIygfo1c1ffnKibFk71YKzX6oQnwTbseE0Xivp757P1h5OlkO06My6PoF79UatYSWpmLFNwZeO
+W2y7NOVC6lrDYqX+dKR+LZ8Ytn4wGOcum9CP19/YT00LgA3tJAHr4k/Z2vtq90fROwNA/5Qo5qn
3ksEQCwwgl5mN5+RfU11sLCRChpl9Q4w8yRRxBbcizqPMJXvixdvC/n6ZjHVUu7dw0L6HW2wjFgb
pfU3Pv0AT/H9RRv7dZCtf1AK3HFS1OQjZGdvf/Il3zUfXXO+EP9/mNud5DV7nBWm5BD1i22aZm5V
FbcYi7Nj2wsKXP90N5gP+qfpoe6y3YCticGKlcr3zHu6jtXfCq1WyL0Vcqov9yQWNraANOrge9vL
mQUCat5nUs+K6IvHSm/x9j1xjGJEpk8/VNEdyo1Q+yh+Doq5HxonvfZoBWySIGaeaAAxoXc1uf8f
g01EwdHomx+XBGtPMjZimJQK+v4KrTe1F938tdZksnS8AKHaXLzAaZDJbXLrjj0YRRzzZlryWX0J
llQHJaT4wPAsGtYA4aCWPhtvgaOXc8V7QH92TSl4hX7nTiOdw1cBEp7fuijdX0O7QIs/hesguWDs
YvpwGLw6yuLZmQMRh6MM/sFLtH//DFmMPJ1dcPiw0oqw6YQkYz6onkIFpNYCZ1qbDcYuFblvc/bK
ouhQ3SxmqF9X/yJeTJkFjeLKAkYOyTNZXsGC7VKrJmI2XOJvKQ0kLTLgzDZ0SIs07ofidO60WgWu
a0n51H6dADjRfSuWF6e01SReVTxRUbn0I2zcWDdXW7aiFmFVYtqsH7SnFiaVyzgkcuY0zt+bowbs
1CzKByHKz04+Iw/aXUDROypDT8nWaKwp7zkFq8qZ2VewIDpVg0xOwnXYZZBfNYKbFGtil+clVxPv
kA7AkAiGtj1o4hqoB0fZ1Y1Dj2rQ8ZFy6Isjt1aivk1rzJ1szpqA9qxHqvLteVFxHS/vsHxZgdGA
UanTvKmF2jBSJ1+H5LJAvrRdrQ5RMuccsJFvdTTquWG6kRzYQYpeDZPl3Avws+LbfcVrJfOgR9gT
xvkXLutUJiB5fwCT6CPHBJrMGwqKs/nz7A+ssyPsTiCooY4LT1wvV1LmiRd4HjNsVetYRt99FbTn
CkC96gZxmBPqeyDK+fr+ZBUEtUD6E0piOUM90Q4Q/rby2FjvkRUYuz9qNn9t8BfgxfNNDlPDjtpV
+JlKxRw1rnwgq+vweq10RfQ8SHl56tnjRSwKYFiMwZ0UBsz41IhyZ6AnHJhDIe5KgtWRu1ndBtAh
9/zS75FjMd4PDD46ZpQD8PpBOEQZK4YSOEwLwvQ70iYLzQwv82Xd33pJWwqo+DWg3syKby9IKUln
dTR93Oesv63qkZkwzljq3DXRQvffqZ6PxkXGeTrFlYHtSi5BX/n/WZR8psX0GvIN9WwNyyrFo4Um
t1gBs7TL08A23fSBYwjG7L8qS5iawjYzBXi4f9xSwRxJrVrrb0jyHBe0aAhoA+rTKdb8PyeKDLXU
9kvTQ3nhPH8MS34X7iPWHSH15WDQxCAP/ZMac8z245APKuaPNpYh0YgOkuzrrb9VdqNlsjeBrcY/
l0MA/LYZJwLNCz0vBqYsaOymGhl/oqJ6NVQxqX9rsxVNatdz7m3MKgBHG9MpQlSHPFX1S4bj2QXJ
j6h2m23muajEBJLga6izLh5dcArxArgKgIUGqZVOO9kALNON8+SmWxhRulR7rQrq6b6AcMX60uUT
KbjszZkwtULsRpSl00x8VEtm8Cl9vyJpsLVXsABlXqitUOXjxs2TY4dc7RjX+pDOu7UggKP2p4d4
VuB1NzrFVlwxX3jB0d6AijsLVslGMVuF/vOypRIIEkApqHiLj+Sk9MxbqztT3y/Apbu4Zbvg2M4a
/vcNIM2TKjCFZJlDBnJMCGNVuLLucynOupj1NlNmhb59VE08F+uFpmPeuiwTzmVSVOiGCXxlOSfN
2KfYFqq4KNauW1UI6lZp9zonPr0CY/u2EzSb0l3zDrOvEcTKnh24q+07nGqrYJPavyW+wOAgV5+U
nT7eWQLXI+7r+G123k1vvmsL1YRSHfVdwNAdrIc8Cj+dxwfTEm0WrSzYV1jAuh68igzpR6vqjVbP
k9Se7oHN0Zogm7+RiuTIfvNVOPhz3MBvTFCaQi5pqKZvhWWVygNTz5pGFz/TufMvonPYGAl7kVU+
2FDqwh37fMaQO0xnaxhZw9zutiMydYF2j06/0qCtnDdwVHj7I85PlDmzuqZdoq95L1115gYoY6vP
P+fuuEmyF1oQ6jzOxzb/VOh71EdGJlB2Y2waRcPRtuhddxD8abm5YQ1ny0OoMTz2a/7O6aGGul9Y
renfJq2hC07/pYgM70dSvVO8XAEcLeF8tp34rfj1Rt4De9TlLITDpP8HCkew9DtVsycnTcDhE/As
LiP1qgjLdVxxJ1Xu81000k2tbwNRUpnDqxhn6sNAAQ6wP99WXY7eT2V7q/a5TgUg1pamqTavLb8h
wPh/YRn8dVlJLWLgqAF73VMM9Pht+Gn86sjvCVJR7E6IuRQ5PYdx8Itd/WeLPFXeg9/7EmceLhk5
KIIfhPXl1HWVDWMhLVyw0EdKBbfnqI/O3JfV4NmfUkuaP2GdYhf5Qj2iq98KUugyli7oXbIRWCGH
ba5wDVDxJyQKEXfBcxD8MqaXdDjlwxiFd8tXeWeNzbFR/OXadYLH1SvPJ/E8EBze7iHGoEXkOdTN
Ek02sw2/tSa0T7p5ZoiudkP5MO3uX1OJx0hexJxUIUHRWyisNbZKVBnsgZDO5QeLM8BF5JUKLrw9
4QPdsJRLJOYaMNohMaLcc7oqsZCgMGbeTRV0CfFlxJFQdBc1NJx4FHRwYt6TOw0ViiuC1ueUgb72
gxYBxgMeR5sAe5s30khGplt/odNXPqQc8eyYj6ly9BFTg7YB78FSoCjZXf4H2xDDQr1+Nlk4VbpK
NdJMOUOpumDk8mQKgimg79BjLMfcLpqSDbfSncZjiMIr5Qv6wQu+c/B9+4/afD09yTwZSm6BjpKU
Ia9U7CgqpdTiFC7uXjMXS81hx3PTAwdW8ay4OLwHOm9NESnUD/LwLY/fuQ7SqgNlRd6Zsc1FW9Wi
4Nuy4ACMRz6WZNX/4yKud0sk0OufLyCX9hv9Hh5KTaFgFeoSM3v5ns80Zbanp5vCGPGxFizm29wX
c9ZIzt/G5KsTgRBIOuewuJgLXMb6U0SlPXhrNdMpSWvYidmgLc98tfwDoSt8jiIsEsdSfEJzy6e2
OakMDQfVjRfAig27lvm92IEPGeDTnkFTEjDBlDjY5bcAm2kx+PNnAbKE1zlj/iFZ9qLsQLt9rJsK
maa4Zl7XNED62DLLb5CKlpnyAUlEUjmAQc7BNHqNWQnrsrJczIfvSkLBrYzBwE5FDA5QlC421chx
1RocTqP8gc214ksmKBftfe13x70vczE2OgSOSzECMpqjgDfpBBJPMd+Fb4TZoIoWZVjDCimgXyXY
PzBgV5gGND1IprMx49WvdW375bMYsXZG1Mh/U9O/spaxf4BR3mGg6Au9eLcB/qPkvLbIfWcW9Ngv
emX4WiOHfXG+Q7F3KVbKx1XO6UK59id4ql5vv7VxVZ4VKu4fjucYFBpmbRsIMMgBajZ6TKXfowHE
qjPXIWvXKpx+FTGpHH9AZbmRakkZboyn+CaVSARCUEggOEWPVLRAYlwTVtytwB6PsR9wnuH2hGaL
zaBDEeNeEcSz64+pWpjIXxlGtBWY4pcMokv9WaEpnlCG4ag0Pkox89EMr/jbf7FbR2I0OYFlMuZu
K74sZYyaxY5f3/fMDws4VN0+XZV1/Hl3PEK+YlnA9Thy+3NePYHhPhWvkQ2MpiS+W6tmxxB/eIUd
5jcLn4W5L4O7x94KpEIGZtdarTsMdIWGYuGsgBJpG6kDLEjEBHuoLLmCv8NOwQVb8Bg6p6Sz/ZL8
FhGZCojVfmdil0XE5GzU5lavKKZfHhL8nfo6hqkkySMZmYPGC8gccD+iE8+hUKxd3KGsE9JY45zl
3ppLJhv4M3VUJT7xRwIk11q3gTmU0M0sknpFXmWgWuyWuUproqVmKV9u1J2904MFtTM8oLR0Sjpn
D40Vot2GB7PTYy0ZdeqnttkvtICoRx75UYRLW2MjAynxr+m5HZj9Jog61UKkY32vo9RZPaaSlzk2
vu40B6cjf3lpTfD0SoEZ3so5e/mkg/M3XQwq/dPAGz0U5O/t7FFNlDQ4CpBQUv3GBX83ZaY0ioPl
Ft5NcsD39HRnMrlGeAEv/tyNaKGppLjBCmJimXw4UuAdGZ8Uza6EXUEnyNTleOUG3cEMKKIr1p7i
IWvdxBmtkUAAOOuWotPrl/NQUwyYS88NZaAd0SQ+bposEqT7MPSR+gJL0h+JQEKRKrV9/izn1a5X
E4Vc/VPPEMMcf0Ciblbq4E5pa2yhyhhR0FN5KCAoqp5C21pSjwr7Hqtv5ZasaZP591FUwbiD6TbZ
xD2ktqIoLNnqvMQJgo8nM+vuF3+tiE+Bz4iVsgzM6hL3WeNaQ6sPbfxLxNxlKxZU2LKteIHDN6p9
TVtlExgEQ8mwRwFlk6c0QgCrwIfYRtdAGnz3LhLGFrrY9af4wHIYzGqAECXqfnaGM0xER5uV6uNY
Iy2qkshzCD+mRGcpiVKY5w3Vkeb0RIJhVuwfHBSYGNkJ3leRGng9SnFDsBpe5tcK5km5NFQKs1Ag
dDftblT8QDgChsq9Xp7c06qD6UHoaEg/ZWPU2aIfxhY04zbzRLulujP9oRsD8p6Fu4XAnreePHLh
skLFBBcS5hYvEl6RupwRvN19EbBz9lkrmQhiQmoaatqErAALD6DguwMmFhIvF7WxMmZIm5V7mPhS
9/qGWa8XB4zB0pdLBZ8JaB35BvnmSJdqHu9CZtm1J7bWbx2F0M7Y2JtLND/pXks0G3o44pmVcjdr
Zq4W5IUnCXzevzhXreJ0cHSASouB0YvjlDQd7zsA+6yMep17RBtH4Wb/+ngCoBxulGCo78QefyBu
1YxPsuCaR5THhwXqgTeaFxq6Sivs90gJRH2DbBH9u+4wzwoObZ/FWMe+SaLF4RQTeNppvU1AnRrY
J48vtVuBFF6Ac0k9xUM1SLfbbf6mnzK4diuB93Pu+sifELzqK7qyW2kgH9Um+Qnfhjp2ZmvLlZsn
q+yaMjF/9RUtUoY3qnmgD184W+UTYzeMBc+g8ij2TxWNkwhEBqghFaq4cdZyFcIbzHCb0ORY9a6x
8COhZUKFcZZff9i5Cd6y18ltnBb6TM9rQ25NWxedVQlnjmSdNWY4xcn3TWHWiA4SX9uTZpZnfbC+
noAHFT3iWJsi587ppWgo0nmgcDoqowdgNs1B48nIzChE8qaTX1WmBvaUWFcVpl8f9j+bNZl5/v+h
xjoJF8tTkagjraiI9MrcKW+u0gUomjODgdombAQdY/gJtCXX/DfXYQnijisto1zJTe8b0LdX5PdY
R6YjxDsf0y6rYOt3PMQ3dtXT44iik9ZjwuBRheNDXxIGjgx048fSm1y/oDTG4AUs/l/8AFkRrIv8
ZWRivODtQStgG2zltgZmOI4YjQSsAyUl0mxQsJ7fql59gA3eTq1Po1wQuVn6hkmSlkUqIh6/yHLa
NXWeHGsLGHxMcA8asPuQmz+7xzM9/l3owl7tzxjiFAdXjPCsG2uJo6D00nVYlj1xo+3gYTh/Dhzj
zxjyzc65axqnknr9KovkItKwqU5UkkEKrIqbObjDSM3562cpAIF4tAYQPUQ2CuOO8+K2zDI0TJxo
K0SHTv1cgx3zf9l2SIvGcsC0NYMRIGybb3laoRpvuIgXKae62Af3qbnfWXk3o96YJNsUZKSDW3Tz
lnIuzGoU496YRp2kSLHJ6+Md75CwTEaRFaOL5CrjxBa/JfTWV4T0llWSWBxchJ4Ln8HkRVzWKBMb
nZtLZkzf4TY1EB4h4VNSnrXabBbKmwcfNwldguAMagdZDiOz1bi5+z1glVd4duorKrzFVM6ehroB
0RniLmzRUAfycLBY5Nh2uAcC7NFeuHSCPtX5DTEoB5vZzZIU8Xgfo5iRySY9LYbpQ42APJInlK0r
5QXv5vzJQwxyGbCNosCof92V0rc8ynyUsz2PYkHpYHZz5PBDo7OF0c4U7/iTavi4C9Djl5EWnUcm
Z3OLk2lg2SKgQSelXnTlgA2YoWhIZM81QjayKDGkM5pbRc5C8QvT10dVn5q4USP2MmLffQl2TAJ4
jeNoTFl+Iq3nZdga/W05Xd0dB/3TPSUB6e6letgJCx6rBr1osnQmN7kluWZ4b0+TjMUhtZ3tgSNu
iifVvuUF9s5a5zDRAsamqFShha91QvHOzPIFmk5pFU0kzxWDJ3dicUsFgoqZbtV3Fd7DVtPHz3Qb
uwx7eGeTDbcMmk+Kyyy35t1x1GVYEYz6upbLg99JVwGz/gAQKjzgtUZGRJ6QYi9SdGPGFC1ROp4u
KGBAokLyfJ1qWfAqHW5GNj+lSiXKmbwGuwyu99I30Jnft0eR0hsH+HSLKE4YoD0ndYn9o3XXCMep
j8lP2VPwoepzkrkxSi63ADhzYwn4uS/qHTv2VFefs3/rVVpMyeib57zVTQibmKlgolt0D0Mlr+dx
GurGF+/DkCGGQ9DpVFOlJc83dxwrG/DSL8bHCksZ+ZNVKsADr1MPGqC1mzSxy7BMXTOX5twlCesK
yh7QChjiYvLwredlYcmk8HYemv4ydQarvIthcpDATgsIqv1RGdmMd14iacBLVwxcLukG0gvb6gb9
5b9lM7QRJ9gKCe3qiXYd2GhmSDRjXw0yvNPCFU84BtkyUzSafsLfs1BHv71lYaHxGOVaJsCTB2Mr
0QavjiAWWtL4ieAZFSyMnsiMlsODW++bhDRgYQvyqrPTm63ZmC0Xc84mYV5AuTu5duNk1u3ztMJ9
Cj0791jQj/KwNvTSzESUEcRDeipBZdo5+8vO+ed5PKkZtbaJ1uiUdqLcFx+btEzpd/c3ELuSJxfA
8F09oempND/xxO+1kGS2jZiAU/PPvr8FPm7fWHvEuc5SBbomUreEbHFXhh2PQd1BTXUMOgjojBkE
3S9v0jw8LfvcnBzs6EfHRKJFVV9csCGkuF26CpcZ8IoRVsbZbg5GpncsWPppaXbDYq70zJStg5Uf
EVGwcTpSHYQTCH1tES4MSjFS3+fg37rttdeRV/HhHsJrLUB8a9vibxM1xTvpW6Vd1U3yMCwDn+CD
0OFAi03q2NvDjadHPm6nY00oNyVNehI1cdUrotiJzFvURu2lUE6wPCY+s2MYe4oC520UJApIx+ud
diicMwUzr5Rj87ODsOmaEZAMubccuCxTyx7L1owqYkwmMZT9rePm4WU5t6bgePkX/gNsq9XLnSWX
kZPFTmAD2xOlCwbK08sHAfd3dtnsfE6qVgZWjNr7laX38bf7E6AtukcVIPODKM5nwxIip/aL6WBT
IzQ2Abph8PaevTtiI9jQCBGHA6kHb5bzmYUYyPBaeuXDean1kgYeJFBF86PTI5ctkzqoeJkreyq8
aYyjjNBqoHsmIqj+Am/GG0gOcQNSd7cLTy5eoH603XYLpKqLYSEO4OpkyzfFtbxYKOQI+MzQXj2A
bMqoZ8Ie8/90EdZLk1nEI80OlSiiOQp7pCz9BXgmf3ShKN6Qh59C5NIwlchF9SQTX2MiAQdi8MDq
I1CpgeLs0+Hh1fQzwdR2+jiiiRXQjQzrW6zsMgA1iZQK9ARQtgoMId/Yd3dDZ9uYmNHUMgNwBLcM
K8Z40Uqdb0L87JpMDnD/ViTQfVy4HenS1IZFS2uTUaf9lRKeJ2COiVJzvb5KtmOeOWwQFdVUooou
ZRSR6TpZ5oHDfIAUztikfRUnUd6KJg0qsY8YaalBICvC4b/u3dDWe7r/AYJSbdcC/FEWcbeB3LNI
FBWqbny+owLNZQgSgrCewiMZwiRNTof8ZACH1hFGK9RnLniV0KvCWUe8Zn/2XmI5a6LrSxzKxEKx
LNpT8cSQw3POw75T6iq+P6ItFigRRNLn1aNdHJudlFOSbVn2C4YjJ6HjBFzHG7aE1Wjbn69Qktmp
7E5DKG/2CPZbge7qJRm1RHr4Rc9C1CqwIfDmL68VLME2iO1TZAkMBXudCiOGvIcapamdC4x14IkR
ExuBSisJKACdwZrCaD3xDitP2DLnCRICBOIbsYAuvkKpNjV0qoUsaqNr+XCv2Q9EyEIBns1kdgMR
Be5F1sRhAaoIaOSvitDzDLGFJ2gFaekmzsa7xuY9lyP5RYVNRAlv4iWAmWd+Y0R2QG/J0Ls6Ko8Z
sEn0K3U22U38xzKAsxnLXlKdvMSl/9SCYOIiLXCxhghNEiqJkAEcfzVOPvDfi16K23hmeioQnd4z
5uxTJCiCVl6TRm3d6RO+ix8nMPdH0GqSfozzchsf/wSXm6kLwvecZtcBSREAt0txKbopKZS3YgJt
4vuW+SJpoAMs36qUObRM43INrZvko1VNjCuLwxc8RI5zF+VHRVOvt7Loh8m+QILsd5gn2Yfkj13O
uTkUETwQoDMSYAyfDg2kg5nnjWKUwyfCSfBIz8O7EMG9h1iL6tHJtahiq7OjbvwxH5lHTWh+toA4
OD/1hGuFs6sYPi/l+2due9WZ9cA+C9HhzBlIsnUJ2UerbucN4umdIOP1PyCj0M7Outuy0/06Vuln
yJ8Mi6XiZMLkrj4ZSAmgp9nQpgOb1rGm7CbyJjiyufu9vzxpOvit4nNYw2PTsiHvPRJI4HgsQBYT
ezktv87SioRPTUl9kT082ZB3/XayXyTxXeaMn4SmMYVWpqjIywpNZQ8iMWOkmkuzyoJW53UAvghB
VZ44UBYU+0fjosa1B5V/s64gom/mFKmp5/52Rql/IQEcWMMJXJrdhAa1VzrnDn7ryD0c+ggYShpM
NIiVkepmlURSbUY+q+Zw98HvnGZWu7IpWPqFXyX6Gw/UntmUTSZrbO6dnIk9Lc1ISZn1WIzVJ+I1
wH9f8jUX+17UXVZcwoAR1BuMVQaBhfB6znRIIDd9Psx4nS6Pk0z7e+yWZcOssOuIy/3ale4mRodN
NCRvj9ZdM/MMTNjODMONdFFDC6Lg1ORyqJl1gCB6IYw9qmsElt39vU7v7zQd+IZiIdn4ZCUfSv3D
wNLUyB5fuDm7phcIoAjJiP5qLkAGaMXJCeC8UtQN+wd/HRVyIZ7gx2juvyBdHEoiRW79haYMc5Oq
gXkIfBn7XRagWWBqfeW6fblLxu7cCP1ZV56w6tAufiLZ5A/Qx+INhEQO5IO9Vbj4RmeuDm53hAXr
dNv5NoDJFrfSEG1vPODC6YT9DXa+p6roh/CMigK1X4u43MbIb6NUcMDfVvwxTE4+kh8KkhSqirj1
ylSlWCD2z67tVyDSBJnI37xfiZB4KDe5FlnS+Ewdq5TJTG5r0uZsRaZt91QZc2cQX5pBvhfAheLL
Xwjt8h1bJ9orpRyahOF4UZ7EVfX8bqEYikR17GpizMUxdAWkiDrhUiTAt6+eSlK8R1nTL0MI1eWd
+SwQ5ajdvPqYvHEucokC6nsMBx8/eXD2GFAIJMmsT+/Y3SjagxP/wk2JYMj4UvNcjlo4QTs/Ekp3
PMycAtV90MStWqGzPcEBazaRyZ3AutEMejqWNOrkHALVWl1DHoGxTNMgNP74LzQ6pF1yicA3KYVO
FiVZaNrU5INbUaD2jAEcC/S6gXYwD0w236OzDjugpjEi/4/bg+lnk3zZtAkV2eqGuLxSTlNUaN/h
pVHeZs1aK5Mh3EAyNzonaB7fzUNRtD4Se1hb0r9ZFal+BbBQCy0JswZtst/oCFdAUK4vXDLYJjSA
Z6oh1X+1T8sgfnx/rtrt63Gm9usGyQNJWtTG4oLyGM4ReAv5h7/XWTvYbdartsUolJbbooGeTJTx
uLI6VWb7wFmi0mjc5jNC/+GUnioyA589jP/qftxo/Q6Lp2WeI3sYMPF7yNNGgogEtlDKgMsJIK8b
mYGT6u8kAwQu6YzR5Zub68Uwdwcvz6jVRsMCIlL2zjvl2EVC84VWogI3n1ehjSSWQE/GgsUMu2DC
69UGn7QhUyW8M6zR8FXPySM8KEAqyRfJpoX1G/ZHl4O0wodw/fzLq6ezFub9qK+rdK0R6l3Qhjcd
eakuapOor5/7/Z7g1f/IQ3LKjXifNKQ86FvEIxqyPVYJhtAMb5uKm1cUsHfjwutqJJjRgczanvZA
GXalJuAouUBy/LGCxU4xH86pN3bPiBfLTAXxWsQtHFa36/lbTr/+l1S5w3cYg1Er+wCvgocRBVIj
gXEqLt5PTOKKVbvR3IZRioPpjnbdnKY60lBtYi2UtY4x4vWkmqkoyRlmMqro3o+xL64l8DIwY4di
v3c/rxvtYJZoMhzDMvfEjpqlnpAvMfE7W7zwsyPCtjwGOfRqmsfKaIx4csldrg1rR4ymosgFqqVt
Pw6cPh1JyahyI6XLV8Kn3F66MWmTjIQfrY6/6VIN85f9NINgC+E8S97KQzTquiTY79Z8QNj60Hm1
ON0gt+HnodI0NMbLEKu8qmhNTTVZxJRpXXaLWTh5vXhaO8GWXO0fx9OTqP4W1MA4qhhVxzY4GL0A
3B83HR1Le61xQ2QYgTTq3AqY0FnpWsHGAOonfxCY5uIfD/Jc7ZGNC+RXPNUV29Kq3xaUrVa0Yim2
Pxf1EqQog6gX6uzYfmQKphGp5xjQhO76vkKWfn5BtAW/WYpShy+plI2ldjplRSR7ZmstMl0AKOyV
V/G9mhYzGRrGwjquQRbMRXGTkus9uTK3mkzhJQVUNJhWzNZ/A8aQBfJpqdJvt8rV73qh07vD6ysc
Q3kgu+6aRJLbWs2whguk3YFPhQXNtORdVt7NwBDC8lmDX+vT2fMZi1vTWLPtRXX6LrIWJMfbdWQR
80uRphTLMjky9sFp8GETIA7DzFhVGmO9vgqHdk2aOAC6LTo7sBIGNneXttyh8OEtet1EXCLAg0Pz
Sc6RlcamwzWbNSxotbK80wrGS4vRnlgarfim67OXKyT1AzkxHDqabEcIIn6Ea9i6Q+/P8WdL2PBp
cX2b8sofH7vAYlH84Rhw39njDGiVbqkHKRf8Fhemks7y9al6UtxpCoBW9nHYq6b31+F8dhib+zs1
PwjpqD6zGdGCb4izdXW4Bl6ls2Yg6kmqibMItWnzByiRw4RrOFM6FSA49DGwFrV5k9PuzgMKMf8P
DeX+aADqd0CKSKTTrna2GLyzseuf54QZTWjT92srPzjewczYas4USWk1oIaiSGEsT9V0hkOesUuG
WVuhZVdBzql/euJ9aMVr0oK5qeJ7HUmEsOT8V2KE9p+nS86N1KklpAO9wEaWrUM/YT4Swe5TL+IJ
YpEY/VOFfsx+gKAzl76UpgR5GkEThqxeBgswOJPseEMi87rrRZVpiuuVt0ZTAG/JFcAFiitVQJYW
QinXWAng9lsEvDQGOezBAn1zXKzRZlDrVA0IX82A9cJKvLnlggjLWpNnKF2GSkM74GL55ghBo5NK
MTOWdcXa7k3ViYH/2SlF+c6W6yCoywfqXjCqkQg/onl1+8wmJEBt2ddsKM1lJjjpEWUBCLSHTOiv
K+yPWvjGU1BO24Yk+QgQOMOUv17xnE8x+u+6ZCOlOHtxeAS3raus3blG4JfdEuV+ex6ByCRuV2kz
vYhUHH/qVrAza/mosLomiVxLAfc5xib1QR4BXuCbSHUpSlwGkqea1zOKLuzC0uDdz2vTMeDxNusB
IBa3UWXQ6q5XZu5sgfGYsQSnXUrXRMKcfFQEOoJ/6InpgXIebpqDa/hHiIXOqf56Td9w3l8ic845
d03RHvidh0bwhc+DkBPfnAp/2VOBCd4mWvpJ9nz4FVHVUGFjXDuMTIYyecRn6AyS87Q3PelcSyeR
Kp9ysvqSghplrtjrzIDjlUtdd9xK1aSmD5uZEnqkyoeEIARtffafYLs4IouqRklLsnZA0+Tzg6Is
qfkf9tMBbc0oEKhFUx5VA0a0v+gU7Upe1i9e7gLw26kpCdgdceiUfNB91HGDMRLNsjvfsyiZU/4j
MKKmy2AfUMnYsoYolLgyrSKGaiOLo+1KkZ/OtTZ6QdQXvaNpt9iz9RDHa/2QwGrpbFoN/6xAMtyG
0vE88AkDZ132ueA8MJ44AtKzXNPUtuf/JFUwlwn9L0eMz5HNt6RO0dptUvmVvyPtDjFCODAndtDB
Ad72AffaKq37Kn0dQP6f74tKxExDXTOoCekf8BpnqmTLqsKqcGilOvI/D9OilHOeobXFgT/pvesY
GxCzH0tHfVLFsrb6hrCrGtgk1y97IaB0UAR/NUqcSGzTD2Rj+8VcoQl12wMIr6Lkm1cq72V0GqZR
aoMddPfI27L1UxqruNYMz8aFSPDRfvwcS5d9qKz1bmIyEIvukTzr7+oVYm7EDYBJqMyr2tATeNJ/
GpKZdxcPzJlvgsojF9sGc6CwDVM+OmnmQzSS4+BC/mBHj+dMY5O20KJWMISXWc96DYePFMCratPp
ntenTjPjsTCuBOnKUT+FE7/iXVASCvVeZAJPWMahD7nYYCjMAnVfq7zI2tFDBTBAJZJz5YFtWaU7
I/os65mNNx4+FaDQwKP3mjBIoa1aeQAtbWpcta8DSL/hhWHODTYMLjTZRzxzUT7k23mWRjOleB6U
gt3ZWNaqnEwjclRJVbhVtfOB7qK7Wq0uW5P7xFQv0coKoMzFYO8ElrNemTwdEcNDhGvpENBxzCzd
3TRhKCUA1FPHzQTPVMhn/05YtfLvpmNQ0rMzC85ZL63iTqE66O7DQnMX2flv5UXjf9AyYztLvlxi
qBtSh054oQVyn9v+bI4WqGknI64KEBqiJthrqYbioIFHY2qkjyvBgu+LXAfkbgjWR/UEvRlzoMU4
gFBary8jfHfvTMGW/JzhsVruJMU58ZRINo5FKbKxrkqVWKvx1YzPk7o/zC0vANDTBr1/2j+hrLLp
BlroTABdxp3UCoDVIQAOPNf6nJwtRm9GKSm8XIWBx76QjLP2zgI8m2BQc4Zb7WPzAHTWIIbzN3D0
WUo3AdfFHUFi+rcThO9Qe5fUvMFr5yyYCZE3wVVy25wCsjhsiR5tjR7VkUsez4H8YkcU3Z8poWNF
9s2cgSnI+rBuPdgUR4ByqkV37cWByJREGIVkNO6iqODyAWparXzrisFoGLWpadj6CQUbsFXFp1KB
48k9oBEsRoJBLTYQVDItde0y4vKosKDB2f2BGM7ytdVDKygmFtUteHSqN/GsQYOOaEGaEMAwPdl3
HFKdJk6Fk0zXXzCD2fdI1IgB6Fu/s6G/kIcWyfJMqeeKEAQYjuL/ihPNJiZN96HdHMkoKrTSVsha
CbpXAPw/hnH9nGpORZ0JasLPI8i+rBkAmxZbfv7DR8y2EIQ8tWa1QqQL21YACGUHCVHN38Fztlq/
iTwuIfOq34ah5M/0pCiAnkmhQyaWjwc6R1L+MmYBVKmX6GIm+iVzENIBmoW10BVLkhZc/jt3/j/B
7Qeso4i0PNNwiF+F2OM/dZf2YL4MplfKdYFY4RnLDK7OEqxRtBh0CS2S1T8u9BbpbK0FpVwj6xn7
ojLxuu6R8kwyQ18HGffdj13SDY2NmiEeQKw/Lbr7WyKfxevgxMz3Bo0UtFlcAO8u7kckqM5CGTJU
yuPWq1BwLs5dQJhXY5r+hK3ZVQbX+XECeA3LsZGhwo4lXya2WTkPABCkYwAHXUbKeC9oz/J3q/c4
cbKh0d/JVNcZBCVBkXeHYgp06pxTnp4UE8RsL2YsnNfHWhFq9Zu/s2Y+2XVmWweH1eJ/oauRt5vJ
NNuc8ieOp1TktY9gdiOYUCFkgf1rclaWBTV9H0QMMvqr9tnEK/6E1zdaAkQVPYYwgU1pfnQ2D3bW
ia+3A6A/89oXVOzTEJ0hwSb40yUZSUoUQn2N2zVPMwCi58uI53zCm/lol7RGDEKBXm9+EW/ziwLB
BbSiQFfhB6p8SaXc2yA3f0BTlxmjbSNoEz/llC0OPrEWLB8NRJXuzZRUjo3H3qGk2vDuNurW5+5i
F3jVr2SD+YF4ISh7X7RRJOw93613QRWKKAcZZKyiXf5BxCwgsOOHMUcJtDWR1WW34lj+OyQLQnsZ
3+H8nAAHxq6CxWeg3Kf0mHqjburhTQBM9Q5rwMHJbmURW/htcbIlrjUV1O+B9TI/DYSfuFb8/qPw
weJlGQiSlGLuY+S1DrhP5dz5eBZVeQIfG5onaiqacEFD+6q+XzBhzP/nJA8RTD6tDGvRkPB55ndb
SN769y8TvwTFgf5zHnLKLRI8XhHzNWyf1pXg6Oq0xZ8sMl1Wq8iukYhx/crL+sM4UApq0SkViYJK
58RhuQ+aQpILi8RnL72lNz0Tir2/oUdm8fSAE+w4lRdjRhoYSBW1aISUDbDjeZ+1kvmmC9yAPEDa
vpDpVje0gDjbcXJtQOqndIt+Piyghti822LYNdpjzZkvH7/cr1Xt7T5qhq/Gqnb5yPyhByCQV2Uy
PRznWf2kTGAUgqZCRsks+XocPuqouXSnrdWCQa23mLOrvl1ViAZTdm2obzDz1OpA3zSLYB9KNe8R
Y5Y91BTN6iuUair98DyxenI0qMxbF0qWu9ok0kdg/vOey1ZsQL4+uZK1Z3j5pm+DM9vD3EF9Fieg
Mz9lVKRb2F/SsUAG22eef2+oLJX/DOv/fuJikV2dI/2NtL5gV6ZEWRZu3vUyi1U2F0l/FiTg+jRR
VzOxy9xyauWYbOqCPyLln8d7/BvM4McZkderDu2OCRk3S5XzVOeICmC7O/NlZ3yiYSfPFvsGMZAr
bbhjkp6Gf7EQETiez2DmU0OMPFPUmiqVNgE8Eh3Md5FGcKdru+FcP33bcl2vMw5oO/O7GX827iEf
fSMexT4stIpR26hZXPRx7hHW9BE/SODSQLpDlrxtfrri3cwM03aVBDpiVSSea0ioJJOqqCaHYsvn
MjQkdcmA+AqHEe2CoFM3ZyYvQMhlIblT15MyLRJycZwOgepDc7gc/TD2z0HPRXRYyH1vce9YSPpZ
lKtXmMawlKd5DmLeeoIQMyBiZwOqH1mjbAZXIScHhz0kDzQqsDcMVQshmdcI0IiKmHNYxJM/Tr25
SbV60+abEypAyxZ16qHwcdpT0e/rVSQYV01y25/rtPDOGfL/klGnex5AyHSbQU2BDWdrfn09pT9O
qUVbFsRd15/nj71Oc+ssyC6Q7SJaa/2qFgtQUP1CGWlvViEKXzvD1BRHEUMJWlCpRVhO74JY8AqQ
7muojA8F69OukscE1HqW4iYSePWDVY5mO+VF8YornJSn5YeWFAU5X37XGl39PkLDuy9cuaKAqQNB
XxMCfExiTRPimUOKj1NoZl84ZmsWhhpIFRbMHp48pirVN1IUX+D6yL6Jj26PmkO7WuO0wSlSm5LM
he8tI1Ae659Gfgx+XMRZBi4kQ6K7ossg8pEWAoEzKqN7NgIAlH1N0jke6HYL/UdoPGzW/mqCnKvn
pc7OoGsT3xG1+sIENESdj8GVRVijQjH0m9vaG50Tp5Hgzwq7NkRqFmwR1TIvvyFJCxJag+Wy3XH/
cDb6/UL9fMRc3YgQlLbwZUTLaIfXwTXZXkrYeclyvoHhtQcpKJVyzieJ75W1bYUYt9zkf3w6yhMe
6oFWHctGIslH50fLaSip+0QKjAswC2LKaddgAgLxSp41IPOYdEwgU5M3gUqwWdCuJ/j6P99NuXPS
t4fGGvYPs5t7qn5I9KGgMSMb8LtrWeHjEf2Q/FfHnW8OgSNmWrse807UvDJLbMnhgZgKLZsWF/wQ
PLqzMeSdQk7BMj2bXPQP5rqn7HJdBbbXaGGfz+BVby4np+4XKhn0V4gAE6MNQbRFPtOdIRPgHmQD
56wsDgRA9n0pCjnFnJgxAAN8ss+5hDX0ftTxMxGri0z0ht/URZMpBlpzaJ/nqi+Cj1zkoHgCjmrH
4OjePD6r7wI5Lv/2PxeBUPsklWMHe0URVOeqfa51aDJAqiJLIdiC6l2PSngjTRgtMkyKkvvY3IzM
k8/VbH3WF0dvGAMFKcEaGKt5tEZtWqyZyWiogt/9aWEq2VaBTb5aPx39DHHlk2Gw2gcA6vmKXSsE
Y426m+rLuvDPObvJaRAVDKZsryO+Gxn2VCxXF3nRL46K4KzHE+n4DSRHHdnOuAmxndFMUmLNg04P
3IuWGNdNB4CWDu7c6mhCOheFAdcT41uguSiIcit6MnXC4DzTEzOU3cmRuRaegW5059b8AchXZH5H
/RaaPFVP3ZdXHm5o9QzhENNvuIsQyoBPTwS+w+FyjawbGuIWAXzVK8pgb//APM/OOncxb8T0IWXp
0aqN6Fa3WTKAzK+KxnVDHwoAlqXu9Zmah6Gj3EyV4WgfoPT+uUL131vNoIFTkwvg52SEYH4s18Al
JsLv1CsMr9Tjzfe1NUPdDNuWp8w1hMhGwFnnRjEFQyHi65Xc6j9/ItJzhpVyessFRCNkROHv7mA+
Vhbfwfc7iKd3330YRE4jt7a9YhSa9W3yChJhF9DxLvhGGkP7yuetF67TKJf+Qgb/3s3zQkubNFBe
MSVv/DVYoqDLAHKdgU9RqtX9/rMYhldmvZ4MXaXBf0F4ShuJ2dIeHLuXufYUr8zJtvnbLDovobJJ
gTghOCWm+2+NI0IjK+Mok50g81FjZor2rSzF4+ObnEFIvOlUeVfR13wB92ph6srkZ2PR4m5X8/0o
qAcoNDDKnL2GgP9uDVSRg9bdjhFisGtK5vce4qaQNwVUYyOH1iKhaYbI+nbMJJLz2SuoTDuqcKLP
Bk56dJNVSj6d+MnZC8hp34V9ZRc54bWOUFzLWxnYDbOV3sljNj8If01Cb3zYo+73koGHD9ZVdEnN
DFKYTOOnQ6bc/Uq2peckIl0zrgl7nxvZJ8JE8NHG/S0nFvPhf4afrrwU5i/h4coyBdR+1z+oSKEh
leTVc8pBjuyqWYGC7lyyMQ17klGvlhvVfjoQzr+3Z8KUTQ9yfvdd9QhB2k/dG3USqdbaEkL7ji2p
lh3IKayZXrZpFgZT2tjLOIJN3cCOkR8qj6X4K/JdHDomqnzELaywoz+3ger/QAc1+T9U8yBB/AdH
4MnUegSbeZdIa2hE+d9dE87/dU8OWnN4NAu+6hENkgmfnezPyOBgp+6NFtIKr7u7thiHgAd3nlMG
WqjG7dAQV39xWX/ND2Y48ZJyb6d+2a1aC5Sv6D3KQI0Dgiwx9EPw8QgDx92Qe3IZCNUvrVSA8TFa
nVYbtdP/t/icTP79TFxWDo/BcLxUlhU7vr6KobbbbXQpFU5D1t6vCFBM3XKwpBa5U5iTYgr+nOki
CstwF26J0+/RdcmvY1NZLddVvI08nb4YvHoonXdxHhhxOSJtWUJM0LqWylAOMNACpt7nQeQf9q/I
CyePiEAUuQda0Gx5SBMzk14J2WX4k6LsK/acAgXJb9iGg08DEzvC7U3BOzM7apZVcJ//Ak54+DaD
09uLdvTbseHfAVasv3/VZ+Cm1xCIOj2CbR4owcUHcSPEgeCEisgOD+qCiUZJcHjvqLVrGTuGCQZg
CUy8/M+ZmgAxwTU+3oOjvI7L3mbV2LO57ZA0ZWDjjEZqWuTN3VhoUpadCojWr8GcJ8MvKTaUplQW
BjCbu3NZFyMaU5YKUSyz3aQNCU6NpDRWHk1yA1UK1Mz7Y1eTrvmNXj9EftQ3E372as/uCPWNoXGT
CG8T2oj5mxP6KEoZJj6RRKlyQrm1ediA36cFs8HTW0akZ8utGf+3cLfrhPRYw4ISjGKym+ngrcNK
XXf3X/h2NgtpaGjji6G+8nwIPc3kVL7JAcS0NOaWpHEyoBTMEM3XgzEqXaLk9t51sgLhDrl6sKA/
BjYJLusa1tcSA2XMS+kEhmbQkVo/9allD441+tm2eb/ozslgvjTeNu8Bw64/ZW0HW4SII3Oh/705
3OkK5HE5iUzQ4zAyxknC876F7HR4jt/DFvkO6M0Ovy3MEwsR2i3id5dciwh8cWAjKWt0XSGADAki
VzFYHI+5uwrqAAoZYSqGF3rzdH05V4EEmRbshZh5qGiG36ttfKvEs6kUBl7aMwcTM0mnFcGPSF1b
FeQz5/LSCuEJTE+rTfanx4+WUypKijaEuDXk6ETS9HQWKcBEjz4cSDF5Dck71w6sqGEJuL6+TprV
kPTVebdUHGGhBmo9jgxekBURR8r2MI/O6sAIl4JA1ITKytQ2k2Y8SjOZJts27nXo5XEwoal83uw+
c3zWOE4F/7/jLdJ3uJQhtRuD8eAyakpWWeb9blWxIbX8jqn+f0dK2VztLwPc1Hkp+KsCS+eHMSgS
DgC4VRYCBSaZqcbLQfIdcsgdbC7lXyPigNq6v7u6UvR/b0MI12qyKo+kcupINxnC/SnDCceSSL8s
ccKZ9kQSB1yWt889tN92n3dPM9camITI8zVNoB3qbpoQcbP3KpMbsiV7plIPjw0lqU8uq7xvj+Y+
NiHbbqnqtnFrYL2CD1PEu0jdOhRbAvELs4dyeJKyn0R/6sv2Nj4fhDPRNix2mEx3102ggPkCuU9+
7scwMcDag1jYNQ57UA1yexkAi9tGE4momOMfBYXRBllXjnmaEhi7+PKiK/rDDDfC98uUbyK3swgr
QSD6FKqETUaZbaIEI78drmkc07NJc5CfaINDk9kot4n94dNMvI1ZrYrDiwiPxONkw3369BO8Tgzb
RY8sE9AyTtUVHSzMR7cTHzu4WNTD6rS8lsCaVcycT4sVcyaJhB6WpN54PPmhN6MBuNbWWP03WEJr
da1uZNQd+/pFhE79uVwe9G+j89+SNkn0ht3s1QMvomwoDJtfngZ63qkZ7+7Y4Wgy9O7Y+E8KeELR
gST02RA01SubD0lE7xz37Zaz1iOH0WqrTuktKzZ9aYgrocJJVft5DwOCTIGa7A/kO2CbHDYH134t
SZwkmhrbNSu7mkkss++IWFVdPbBLKrDQAOow/P7xvHrukCpzNZUb+E8RLGsyEBhYiWUyDQ2JB787
uFcpKvVa9YOB6j0tRVRCn4XuIOfmUoBgJJepuCCR5te+kHeF7/VlUE2XokzvZcprkebzwhsBRCja
1BtIt7j8LBMmc+crAEChbEBJdu+Qugd35ZnP0Sg1n5GzMVcVBrcb8LvRyjBCoqA6BXdM87jyRYJ/
JDnCaSXPlNkQKJ21P3ElJcyoq9IA9S/jBTb0A8H8I1iTAeNqLEUEqWJdo3B+0mtJ/ooGivANh3w4
OGcETNzSUMVM02/42+1D0c3/cXZaK4Rj8izYiLtYlArYV/vKCQR/oJUBa65xsd9OT0nqEHULQhIJ
Xh3d4Qogj3Cttyu0CcCTyQYWbEAaRiqSFGSYzY/D2/3G/fJ1jKH2Hu3mFe4FO38zPNN1A7OdbBPQ
eY5X+zyCO9ii4tOwocxwQOLY7APD31k3iuz1VhYjGUncIZSzXwroAcJaTyxDwMzj0vHtWmOyZj0A
Dqm4Np5Noa7I0a9DP75ZHdm9btu7BykesM+ANfZIfYF7vnBfiogdJLazZxaujqQjoAlojulxSeL0
6P9Kkm7bKg755TWHO1hQv7qLYcqvZ6UVGH6UKEUhrxxvs77BYkABqA5WyuDiSS+IH+AVKoauagYD
U5njrK//E37/DUTto5LgOtRtY6Aab7pkK9RGKOTK8wW3euDwNqN9SqD3o8aNkcnZroadj5GmNsDf
JgipxVoaTcQeJObS4332bQH0oUjCnEpPAjBh8mHJqrTPoyRE4V6IqNdLeBpgLD3DnDVDZVT7vzNQ
GGRkgwW7t8ipzz1IBhSKc6eh0OgRJgJRj/s0LLvkIBQ35yoz60RudWr58zaNRsWSOQK8ty0/rxTH
JoE2zV6Lrqz6tF4Xs7uostMmLkXd/JC789gA3Knagjd4rKx9GDEc3th0KEXJPzeImeXSwxC+pJ2u
Mh7SQi7QQ/rhDPJ0cgPca01Wd0bJVxi3r7f8aaxBQjbHSwdS2lZA8GJAvstTIYNZHZYrhgzzjVyW
sJ8LdDIAQkXj7zLG0uezHLZqGhdAkIdybRSo2myGmesEOUBNnSirB36B1YgL2KFWryH4oVKbln0P
gals5u407AMyMhBB3iU+lcRWSPCKsqk++ClmfvFctqQf4FtZ/SSrDo8BPuo2QDLySApSk9ZbfXaA
pxiF0PTfoz8Z52hLviE33OFcd/vTm9r0lEsKbY3EIvEtT85BHUzuYX+4uJ3UsRBoqXRCGq3FF9U4
/ka31cTolAeU7B1O4GHxHFtkdGjsINadht7Mdb1RN4kDD/ACW8e8iitfr+JIU9DUMvbNO2ibvSLL
sNhv8xSl6+uCHTKWQH39jrVDTNyPyYQWDDWs1XeuaeVovSg2GAOgemDS8mfz17pCC9VN7Abuom5h
Ja22h3ceNwnwQS5Cis/o7t8vrgFVLW9UUqmbe5bYmY+PrVy2pQbBlKeuwCXRhmL3tgiqIpaAMCVp
s4r0FLQYk/d7KrSu+3RB1L08gBwXVEvYXC1YlUVLkxp2jBa0VrjGFxaPBVXE5UAr2tijByvwMqtc
l+4dOlKzP9Z9yap25M2hjgXy09pcSsJXJfGYfRysuqIpJJXPMQZg/OQE8tutNLClKj0WZw/Kwplm
/givpeAkgW7gsYoHJ1rzjoNjSz+cTRysRM1ciIXKURwwXSzLB3fSQdEXcgqfjO9hSOpdiMvjHewZ
4YIl1ZKc90oBaJS11lTwC1R/mF/H7zAqkDLDQ8AD5JpUYrQfJ8zBy2G3+/FNMSFveBcpqRMJW4f3
j+FVfFmuKvk8RjSEHwCSlfkWfLudn6GiZi0VlsZLi08JnR42OqG6fo/ju06nSK4qCooKQ+2D8QFI
fFi8HE0W8L0C7qRGZNcifUggN4o7f2ZOzCSJTpnrldtpAp/Np4cYmGQM7fhqXQzLLmIhz8rdvQVW
rEiOwkp/8s/5k7vLTKHhRpLY7jPnWDw4D/zWAz+qafxf/IBn23jXgtf+wAINbgzmoEoJYn/2e4pp
waePu8Qql6P1GZ5YmZqhAnrvYWQOnP+WoVlyGosUCiq15zE7w4YqoHkhBJ4JJB+jeTJ3ASTqau3H
8ANOTbtWObFZwzMrJZhST5bBpeMF/1y6o6IjzP0LRLLa6wGHEKG84p+i/dcB+iDxuPkRdoC55Nwd
qgkNOSQnbm0TgdFKNM+jRyxOyqjrm9lz0oHovhJzCoKnbrvvQSzXwcCkKa9HDAbJa4XFotf4fuym
zMN8WIei7fefoXDBYE3U8Gb+0/Eaje1/H2aQofwr/TdBB+1AN9AL1Xw5Grurg9RAWC/XEVRj2Hy7
Oqo7Ch+1mqeRb0R7VPGx/bE5T7308sUcIrjmx1I/y5/7bjFFvKkAk2xDfkg6qGO3pKYbU10b5wmr
fMjPfrUb1uv0k+xEVBL3wrZ2FFTlSB8e2q0c7Ra2YuNK3QG2PYGhW+/NPVoGHANniRGeNs1Ee+U9
EKnhFHxs6nM6nLnorTrJDL0vzg3hR55EPgieZOOgoIqhhfEvpXBaDb3wEZerlR62mKr7a6NpQcVa
zPRDvDXSMNOAL0XVWjHocWvgJ7LJQ7gArAmXYfzsE8JHBew6MsliJ0531qfOlsmW9Ya9lvuWMmA2
8OtM6IFQl/NkxjDGQRlJASCuUPwY4zhlm2OqZgcmoeaS+G/CMYcMQdVS3amy0qKQUotWaOmtrYD+
RWsVHsJ80ilUbZhjuisltUliy09+i8/RPmT1CyfpgmFXlY7CKAirbzkOjjjS76ONQk6rE9yF3Gyr
rAK5NdOr52WFSLxqFmla9bpSDzpP8kysYAiQBNsyETtQHMOc4iLtxZr2f8BNjYDCouu5BAmJfpbw
IqXwG9A8uudMkz9JZDUTNVrTl52wrIGPkaaEKLJMHUbePVacrs/s2p+xGjpIaoqae1g2B8oGklVs
YL+sPj2posOvwBfTRmRmJ9U7rt4JmCkLax7mAd/ZKShww8cg4mlnW8A9/rERaNRvLC5jRnVLDPET
rMfsyj4UgPud+nMBSKmsUGHuk3zClEzFM6saiyzpWDEz2ZJ37TyH7aO9asQ0ajkaxylB1IGcEJq0
B00rt24Xy/++fxzd1EIK88rVpXp1ug9kpn6qBchmYPXDceHwC8rabkoLubmTq/VF6a94iIRbTrrZ
UFNvHtMKnUq54TS4ef4meYbDiJD9sv0BNjycLSlqs5Oo8LVletnqGmUGQSQQ1hJ1Jx4jmnZxFkib
W3R7n9SApJmtllhKexIYEhChe7onsA+cIp+nXVxf2uKT1ZQG334JeCWK691ITVPdDXKMbXCA7/vx
vKXSkPREG2KDfHNkkD9qeFxz2pD3hVesQoqVp1bnVfb6wnMGjUoqHLOuo7qg5ZKoPUEnVDDv0+zV
PHMQzJ14qujLB6rsdHY4dimQsohIVHfzvKgxw4qmWOb0IF4hsyh3ah548+3Ceo9y3KD/DAhY6Yn3
gPvbjxmdrGcSVPd2QWEL5pK1ycjDkmFDlw6YxuHe+dTpVOfx+gRAfyfZuJzUF6aP7x5r+3ADMq0s
0R/gF0Vc+TCmMvzzVPSQAdw11jiJBq2hfHRFU+ZU91Y97t4dCN73YkZw89QE6oElCGTew6tQ1PkT
PYFS4xXrhrRJS2ryYOa2hpTFVAfSaDfqjBYgmaFBsYBE2D5tigAFbzZ2Tmz9H7IGR8s4ZviV/ctd
ou0gXryhr2Zw3HsKZPhLOATkZFyIeMwdwVd88VHf4tmRhDW7XdWrZq8/FqADfWUvAq/R9mcsfWOg
RwLPRt3Qa6zYuBHjenK3DjJiwtwHl9VIIIGV7bqak8YHpH8gm3qjirnAJSeYN1/HHQ3ZaL77vFvj
wwBWSw5pyxLkQ2dmWnjYbCTYhnhBNiZszB/1kHxElX8S+ttSZZzO4eB0E8BNKCVhdNPScyGLLZjr
jXDr++f44zSY6JPRxL1liI0AzhGEPcKtazdAUQImENbmwLU7/WOWGl5nIb8uuP424VEzowrJ/0j9
q6lDIjtem+Cxkkca6/YN2/WLWUeg4G0eaX/KY+yoRI4WxYA2hBdTUW90lVcINaKeRAUr6rtOOfN+
PSwM7ZUiAHPLjJdIGYlwcTeo7NvsIIeiSzc70HTthAyVXuXySDvk06J5pVXAxf4LicXkh9FOKnsg
Px+DBznzQPPoLbKyrDQfFcDgiLztFb+g3lcDXldEr0hZcB/rYEhR3hHHe2Xfr//N+93FpXvwDVcQ
iPHFkuucgt+P83ew1ZIJ30iEoFTSAa9qci9AUGPN5wVEvAATGjcfnrZXcG87iTnL5Az2lwMnqrVJ
/Djxfue5rl4CGDl+7wzPr5r5dEQwuVNjl9NVOyaksIckBm9n/ctCpY1+r96MtU/on6S9AF/Jlw9s
YXosuDuawqDpUjzdOeVKnM80pmGSvoF2EO2Ew2wRYaCZB+HlgIyRT5e/xJP+gQ4IdWwq6t25b298
yrwu19JmOqOh6vYQCgcvVg5qr5YfRBjm8dckZ1qLt6QOibxMvfke6ITpn/cIukd1GI4336bxvcEG
RxTGVkaYFDhK+C5FA4PNEtS7AuOp2wXb3BynsV8FbOz1jGoLBz2lbKi7oa17FsnV53+jNfM9aP9t
Xv/3X8ZF/g/9juHRYWYAd59cHjo4lp4HnoTM38CzHiKZ6s8TyET6cnzp0v12JeR5e47rl2TTGT+p
b8ldGxaFxdPyakxxM3/RxYHZXceesLZ5KwuiLF5I5ZXnY66ts1M6H+TnicoJdqGRrWQuu+mlWIjR
Q7l5dma8RLX5i3UmTQCcp/n66OHqFdGqbAYWIHME1ZFvVpPmiUyiOP6vNAD2Wa/SIMO41EbWanH5
IHvRVPW968MZLIJduTNk5oCd90rkb01Ox0+DtjrsdmuP4Zz0lJZkWGoOtvV/SISoa03miWmMFwjp
79XKqpd1fRVIc0/0CgHMzUIEuPRSf81NXgXJaU5NWJC9U8tPTrelcM5RRwwM0WTFcUNvSXCQNTCJ
TUjk+X1JHqedcFcnXPzVrxNYN1tsnESq6rxvpBgeC0x5XFdo0snlkgek5i44UZAL4XM1jOPI824+
d2AJ8ObVStq0xqrN0nJoElM64i12jHgkA8YDKRporuJME1AFPKg2kJJw+pCQRZgrVb7qIye+RxAr
uJMQ4QX2olFYkylpzjEsEPxCP2CWOV5GMAavd9JTarF7iU2EKVI0onIfTMihWEjlyEwMqqXqIXBv
bJ5fmV177PwBDLtiJf1PbOIRp0pAefRPtwpR1bFkxmnqqPLmltPcOSuoatOaZR43csbILlEo2gAW
ckzzy1LgxbPrQekfUQRyVTvUsUj6fOhiXnBxDiTn73y3yYKhv+z8T4GtmuEbSgs8fTzZnIzDU/7H
PHU+UbT9Vtv2+vDa3ux1HE2MHsebqz0Zr+MLYVJmiTlC7peyfrbXfAB9wOzPBt5mnoJqVCIXk5YI
wkcB0sx0P7REV1QTeGTY5JKixw5Sdryt7dYKxQSFJqudEO0bwDb4yxE2icqq6eMwodW/ePEtm1Sx
O5ba7W3MAUJhBo2Y3KH210JO2w8Vr+pAbcRAj9GkOKVYl8YQL7hBSRcGgBDHfksjn9UERidYMlLm
bGHAVflmUnBWA0Wq5uSGP1PYoRhvF/bRGFy3GlrFrtPmWMdjGZe/+f/gLU/GqbSqwRVwoH+MQBt3
+P1SDblubx5BQZ4oWSpEBH2oFmdcIKMzJs2HZKJ4imo3V+ZJ7C9FMRSb435uX8KMfr9Nk7ewq3yW
S2IYLKCy2C8k5Vx3r7l0MnLk0TY8PqNx224m4wukxCsoNMki6CO8ii+DEwaOWpdsDIVYbtF1p1fh
qtOrlhqWmkelPS5I1FRSXjEyB/2sRXMw+T4leWk+PbjJSD9dl94Xe8G8yRUlpZXnLSLPdGjyjH3B
ReujY0PXGyPaw2E2rEdC1gowIsxQgt8nUNnVFtHH3yp3Vf3LTSFORlsGoBZbAaN3qSBivDWqe4Ni
4UvWNWynW24zONp+xl5QktJQsvhqgrcmrzn5zheP3dtbzABOPa+goNk+GlhqdDYg7y6Cfmt62kfq
FjApliU+QbWAVGJFAbNyyIaMnl4BaqIZJstIlv8+5xNbSMAyWhkvetqD3mCmZ+97Jg6dWxFtkKTx
PgupQsFYpWlKZV/nrLZ6SJE6FtPOSZI4fvQGW2ypu/4eh3BGTJXBBkxyVPNW1A5pu+nb8S8F22Ae
oPhpjJnX0RoLRW5m5GVfn8UIBXbaABX2fqvdREf3cogdJwHrDNkezeo3CDooAbkcmfcbPkJKDXf6
DpPA7K5+e55VjuGS0IB9OW+9fMTXVLF0PZ5jxph8PKrXbIMmqatA8b/RQU1ZHsb4ueHg57oUktLl
t11G/qv+f/g+Gd+j90KJ/VZLgOUYQ+dpX1m1d+xNpYB8fBUxrfRvnLjUbrkjjxf/if8iH+OrAuiB
uiDdxGfHhpnUx4zSVJIWqXStQJRoLGxGIYUJmyIb050ss8vMT32tKlCNyCPMBdrmp+F+SSkBPcUJ
6n8Z/WwUKUXLqY29hhWqDeyFZOky2+Lb13DAqG/EwIRWEO+4wKaf6ThaMD9b2Ad/9vygMOlnlL9j
4z1PGHsO75C+VbDPGK9ePalMyAszT0BTD6qRwv5WgLUqW0+SkcJhZYGWRmZoUBZoymqBM7vZZqXU
Y/H8odbVRttlukd+eWzHt3hvvYR8wirZGhiVH234Pt1ahAbyFJ9qEgPL7IANIIZiVPVtWeM4ywQj
OsaqGi/PsOjpjvLjN2U0KMGHTQJb5HfNh+5Lz/uQO9/g4oy0WJbuRw6XfTEZBudaJwTFG3aoDUYS
4o3h+NryazOoAvB0uWa0jREen3Le1gxEceV1i2YtuEc5x2btsqQCsd8jKl2I7R8k7UTraJ5D3w5l
sPQ4dvfnt1UI9JZCD7OXmRC7wSeO14g9FJE+5EiciuCgdlbMLanYQsXWESCrqUNYecFaPz5dlYnY
LhnjyJsMjuK1kbE3iuRqVMdTXShLv5xKxWWobSeoNFe0k2IMbCAB70wQ8xlSn6oLVX31s0T5JIOJ
sivyE2TDhe62pIWUYITN7tJqgkYkxeHoiLmoOouDosgnJnCgO4B5EXRxBdZjInX/gfHbYlhXn6ad
66kyzsyUCVRF2H/v+kyuB2n0GOHKvyjP2EKyHOIvvdpjdRMgLvD1EwQLdbe7qWnWHzAUIySGJJC5
F6O56aVVNbPyhmqb9bC2NYfl++UP4aGUUho88txJWm0IWABQcFCa5a/thNMOMgtCcE5hZHitglQI
1XMIpMEDnoSz4KOah/6gEuvOtQdiFoS2E68C1lDcWdRry27PqKgZLr50lS2o6egDLKe1/CDvXhEb
hJOcA5tFACSvtrvPsBOrxqRhofHXTdOUvZGtovddXQ++RtCurI4Fpq68U0If4kWKOtbcB0SO62Zn
FkPC+QdtEShOuxX2moThCPz9nTwR5HPmcapTtjexKJyGmcrz5h0kKtUwHxKcxEJWsXuK3uBu/QLT
dqQyMmrIdo7jKxijRdUgTVlBgo1iTVxOtxzJ21/i3N0Jx3nSx72Xx3xlzeonGHxeHJ2yQqEmsQAx
JhCHx52IKaJdKXPgQSX9dSUIPl3Yxx83daO7VssrqfMxanl8DcgiR9HpAV+2YAKSMviQEdrDmihw
/vuXrSTqApXJhnTd2WHfPAZWNLwD54WPusqPICRLhf4oE6CFbA8d1id34Isu/GH2gekU5kG6uG/M
mjuU6gsiB4HuLdBLzC9ZlFrZGa+vPbgZCXfMAg8hGz7qU5gBAz9Zz5q7IOE8BoAiWOd3sQYEE4n4
/UV2x1DzdHNfOQj9yVOsXHSx6PlCNWTawipFO8jZG4VgB5zFrXM5tJfTJF03+2bI6/lRmzRt+fT4
UfvzTAtl1Prt5e9xpF3pNeHrDr5SKyB9mS9/JxTJPOW4lBEgmLDsnWju5TpFpyx98tHEvbyYSQMG
A9KjBNVOr28s2SNgG7jeAZdlV5ShhZ2d1cFs08nJpRlfrU+wlk5t9kz4jq7o4O5ulsttFJEuOxK7
ScU0UaJOYuiOPjJLkgeM3Y6ExmQTgH8xyP+mF2t4r2owjzR4Gor6KxzockhP9rLP87j267bL9MrN
lRfiDoONb4AUl6aHRtkpWTlstyDbdmWlXMAMOXI4kjPNSGmw7/a+lH5V6azuAocfg+SdrId2LwyO
ZUZQYCuzJbKtGfzoEkCoAdRk6vldzJCGg/ZQxKyGIBAQ3w+j5Je4+bwskvKSD8aVK2jTP6v6m6+C
58GAYXxr9GjC6uDljaJDTNw+gkoS4/iDgMoCBLWoyWJIZwd5R8NP1WfHc0eI6HEhnL+lFD9fjZfD
hqFiUsGK1UMyGY5Qakog0hc6HuX8dnjZ4ptmn7vYkywDQI29x7P+kJcK5OmlE/HdQum5h7GgNYYB
CqXGZQy6zhxYwDNfCJz5yYgplARN6+/ElxPDPiKh9QQiztomf8DSfyVFgBN3lI1hmUcDZjucrrMW
ai59NAccvlH874m4hSh/XZIcI3+RKY0nTPPaTP7WOpVS8YLrcTsT0wqGoP/Wd0TPa+qk2ZStoaTa
F8SXltSJzEQ+I50Mxi2XvNQwiVotvqtAVQldteGZQqzn6Gr3ooR1JY8v3YHuyepCHtC2IYJVWeeS
7hPSpfq/qcKayU3Zcu4MjUqgyo50uvRMNJgJqvHWkm0O6lVMeg9NNwMeLhlHG7g0837nPWvx3pP7
gOG+I//6XJF+BN8EzFySwN53Ed7clCbyfrK8UHlo2UWIuMzyoBxGWqo+46NoIO0hm2ag7SnzRt8U
ShXI7k+3CUQwW97W+SN5z4qTNTeBlVSw0hHp+d+Be0S3aa/zJns9RX6KPsc0AKgXYlIV4E2ZC5Xd
KyBFr1U+O1/aZNzazC7i2ETijOmmmILOHoF6InXboGRLpIy+VTZ9p3BtJpS8yrAEncg/GmKKQ+Ws
FLE3nIP38QAQvWL/TAG/T7mqNTL43kIAiLK4FhYMu/iMNkpYTp1xjhi2MVwbkf2vLDQG2XwCGEOn
yWrGpqm8QtvcjIP3lz++59yRKvf1F+DnveF92m5ffqiOnhmZNxQEyZ/u99IcYkuiywjl1Fb5Cvgo
3mFyuvpBZkQRtQxyDzk280426sf5imnGfllFaACAAlW9KBZ+XBV62HzZQ/EQo1brhtZxACphr6/9
jZbtsR3lP6nfTpVayl9UuCfC6/fZUESBd7kT/+QC1E+W+avf38kBlle+n2hUTSbhflSckZ31x9GI
oI9guroGxTnJ5EkDjqtufaNQB/teMPrtkgG5CIlvGaYWFfSFaEkffVbZ/PCyXd7+Hc6vqtAHSN1n
jck5q7D7/D0vYnrodw3hI9hdM6NtPucfjiyx7ORN/Zs79jajrrubBo03FQT0I2qVMz8tPyfQFt3j
GRUsyfpn4JI3W/DszE4J49iH9ER8khuAfnoq8CT5fKwNTb1tWvDZR8jYFF1HxPk5RYLohAja4Ub6
lCsexvL6YFmlo3NpSrxwGV3ldYEXcb5Oh4T1KyfucIFMPRtgqvIuF/sTHCbohVg2F6NdtoRXh+vN
F+vORKBtj0+6hzNc6Zi8pkccwi0w/IU37q4XCODp7bGHyxOlXqU3Bn2c793QdWbBU2M8Ne3mFCP5
HDJSDdRrMzBzBDuo04p/RTbeUd7UhLVHOj0wlkw7MpwSY8sZDYv5eoDKv3VEUCzSYlQdNtLYDTK9
8YIm6lF4P7cxGICn2We55RU3efxW05rP58yETdIB9qPraoKmEL2it77XlMBRdtlBTjWInmSLGzwt
ufD9WZ3EDuQFebD/YrpDO65PHhsrOMR812hH5Y5go4FVEekc8JzB/RBuLtpCT9PvDqLn7LGSps6J
At+0p3oUvbayoLy+u3Bdrh5v+Udl5TT0BLyuUSdNpuT4XIxoSWb6VhIYigIXGOsoMc6JzrsVVrxW
0N6j2bPj31aZD6nuZeRLNddStqoQJ31NQ1TYUzamd3ljSK4fMDEQcpfXqrVYPLRCxaeIsE3o4RSL
VveEySJYdoOmMAyLez+yupjKjwrd2R9FE7RUhWQoBzn+lR5EBeL0xB3ywK661pOff743YrUwakOv
l0YY7eJiTsEqHjY9DrPA/pagrjYLFlxwarr7WgUAaeYLwVQgJ8rntwEgz3TlXKWQcwFmqHUNayWY
N4lNMxIFT0ILZzliOZLfpV6vlIE74QaBbOUdcIsx7ApZGzmBsTpr34kaeM9mlqOkZXV2vwPLRnLS
62DIRowXy+cP+DR2djPl4w4h96CIKjJ0e+s5FfUb0BtUb4sixNa0z1XAfmw2Oq1pJB/r4hj3xNIJ
NCEKYiEFqdIvYyRD7xg61w4v4ju8h6npdUqnySUDk/UbTMd8OarvqpcadAEnOLxIqhRpWgYsxWmY
QjerOu5shY7uvKmjXMncdSrxMVJyKBs9iPUr1m7oYCps0TqfkYuG/6NGNZuj0SjMVfww7J2UWUlm
t7JC+9zKKs9bahrAEc+qnpr3PT/R5RmSAERB4pA28J09zozRK+IvrhgAi/84CMIjtlGCoSPggvmT
YXCpG+kPjj+oECV2jgmYVr8VcqrMNyg2y93BJEszfTj/Paw6PgOsgsLYTHBMs7EXHr3HHnNZzB4z
an6RMoi/HHdvFRpeN4XvrOhKlnnWxoVvPWpo0FpTxK5vLfDwsxnuhhhS47nb6rIa4L0Cz0tUM/8g
fZKATo6uI9uBd+OnauwrBbwYoocAEFGEaGWyJyRDfFbHhlvbClFxaKGCrXcGz+3YxflaYeThzeEh
d5sHZqCrVfdh6nK0lVy0/kYVNrf3WbQi4SzPPF3kL+4CtYXyruabkBZk9rsWHRMlULIcN+25qU0e
+vRIeA4Lc9ihVWIMu1WdpcdEV7krK6yk8eRRNONJ/454cJ/ViAz6qHvDr7vdMw8KVofISovtazaU
H6/Wqpi1J3EHgzZjMMditvk5DnEhWOn2UK+286BXjS9VxG8hl1ebAdw5HKt6ZobvsJIuceDwpKRw
/OjXfmS5M3BsQlM3Mt0WPr3mHz0JnY9fIj3OIMrDo5r9XtiOWAivorp/Z8tTWCzzTYik/K/FJefo
VNTzXbdTME1Ofs2nRXBeBxP4HIEK8ihpNUyrKR2RZnSpAYY7+W1n9SzK3cusuQ4BrOvjdGU2s7Yt
tlb3bHefsTlfwifaelUwtNY7BRJu05YFKmfE3aVgbpCA8VgVoQHoCEP5CYGiAimNpuGcKmRNmhSL
oErqw712ilK4eX+oOdQ8xlUers+pBpprlg+D6zgCovakXGgfB+9PDFTLQUCYGNcDgKbdVghgW443
RnerDUHLff7v4RdTmTf2jJAp27iiCTZTYiBmFJM1pG+QjCH42vfOJjHCG4gi/NY1CUaY5fg75s6E
Ve1NmeSY90CDKasMhG0cQiiIG3hzIjXcrADEJW4aLKjPEHoLKCRHtT1DkCAXcvTwH0mMeOxGYtWD
z5PhTpzcMl9IvVy4jZkc65xstb+LTl+jqnfW1Ybq1yu4bTM680ceu2Ae0nBZx3PirqPpLZUy0zrr
tBqui8bye+xrMjPZ2O50ylbVvdNt7SwCpnzHzTDrTzIv52M2hT0mdZI2T3p8VX65FDH5k7sgvVLc
2N5CeB+PqT38XvVPjFI9PSi+1LtCU1GGSRnGZrkMayTYrRpNWXwPs42CiyyQRrTTBEp9gFvaLJBR
A71XGksxslXGXnQ4UpiMP696qHlc2ZA+htai8CoN+w+xy6IBDNGkA1kX0fHdmHEGgOeMAE3a/rGw
1hZQFQ7ekUBiiGsJgRBHscMFkXQH8I39td/Me8hOUIDhh4N0mhO472KJ2BXyCO6wuN0VsDrlrAmZ
ezltt3BzCUA6Vzrms1Vq77nEY5QRFS4iipLhOP77PD2bqwgh3qkgD29HmtXv4vjxWsmHxNKnUJZN
WSK0Ly/qSP/lg6Co66mMHAIlqG6ZEK97LkotQagYRso8HIm2aT8DFwQ9gvNZmeNBhvH/Qwdl5BjW
E97tsmtScwRIvTEmMAGBOREA707YnPNO6ncW/gMy7PxOiJoTpTqDrzgHPZtoduwXvwN8bs4uiSn3
8oAp4rE9QISWI3WLoUM3OXiZ/HVxnwIteUTeVzczkjdPp/jIlFmVFwf7wENTvLb1+RivT7uCoOIE
cw/PKeenTpaWZqKtPvWTJ+97PrBX/xQwWMdqomdxxyJj8mM7AmNa5o9Jru4ZFNY8T8cpAdxcxUvn
2zYYLd8SOuZxBRJYTqHa1onp3rUV7MSDdqKrVdxHzWC5ah/NmXLEGnKtoXh5Sq9AN6U4MxdAUU6R
EYSt5uYyJlNmWYm1f1TmVYEXmeCMCDOfYNGZ+pKTxtEBl5OxgQLQIRPy4/bJNnSvb0L44NjP7gqB
IkYrr7RQ7UNHiTbH191/cHaQGy6xXG9yjSLSh321QqSUXc9WRAOvPnEd0HRq7zEdG3BLdWHxhkNS
vZ/omyM/amWI9/J29vEL2Zdh9VFZodcvtqQ6IsGUmrw+srUeMDEiZgjLiweVdDHhVkf1iZ76qDZ9
p6kGjMwVfxH6NnfdLuB0LHaNGnezJedtBYGhtS65Bf5VU7wlEAknwqUaAuKwRuAovmD74tew3mC2
emhh7U8Hw3lgtPPCK/kSYcLhbz6GIApwNFO8roVvsq0kMHwPbzT5k1PFh3r8L6Tq9kLj3b6YvlEr
BxUCFtyAAwyzzsBProDJlcuKV/j32TEMMuo0NdZwyuhMTZ8SjGegKqa/A7pALW7C7x6raOJUMeQa
Kw40ARLqiklHz4vWBSfvrsAYvrp0dEKhJhHVF3zTVHp7P7r/mkReuqNhc3cH82B5jxlWDpviQF54
DgXEuojpzF1uHWXzkocxZpD5HQiFs0ilwS8L+0cMI776WZsiT53yLhU5HAoSDkMwyYTMQhcrpYv1
QnkOMtqcZyhug7heu2URdd/eH+uTUfOa+rgRQICgheticHvn6ks9h0wvHAqNmu1hWpzyPxGQd+ex
nqWiFOwyxfLi/5NeOE39tb+keIGRj1/Hfoss1VH5LcFTCE0sTZJ9MbHtpV5GIoulA7DG1EdUoM6B
MMYUQSyf72F1Rjuq1j1fjgS3EUD0/riG2pZDQP1aigrM90zQ0Rbynw1KDfaF9ztsb0p0HGwwt3jc
6tSNd8/124zvzmak4rMv0JQuFJHP9j2a2VJWMQB6uiKChcQyQsxR2GmskDKgA5X96ettFRHVzMB+
hcqDW7gV71Xmps7INuu4RKsJZIx+qVhPFjLlWeebE+mJ7uIyqw+vRflLiBpocaoQuEYaHMDrGCNc
MzrPc63g8QCU7OY0W+lhPV8aWVzMqjsmcUZv+HWS7NS9rdUhlHOFDViwEPEx0xnzqMdMHGraSIVg
WyYtc8i6VVsLRPaANBoTamYrK8B/mO0f0C3L16yybo8q5DPJqO12KODilhUIao7OsJUJ+00dUJme
zKEA1gsuOrec/WY3N3OFbaEXcLiRbRFFFSJpuKcjkk8F880xxBlulkSMprgPQsfJZ14XIZqLL9y2
9s4v6dkvkPRx2pOsgyOzQZcf2O4z9oZjzIuNZgqJYydVt2yz32dGYorpX5g+24LvyAhSj2GOXagF
n1yMrQg2O1wrBPS+TXrEH0buCH4IiJ8bj8L5nI2xM3W7vSZmAczLBysKaPD9CASBkrG6Fcn9oDVA
QuBu3VU4TpXi09A9DYTBv6dD3GGFFfeMU6OtmyZCoXB/+3rbE8Rg0uZkqj318LW9GBcS1GV4Srd1
LjYSoC9Mx1gcsKc2EGE2E+ZGoseGcFfqtBxVygBFg9KgesSQ55smaUTenVmGDU+5tMDfQH+5kwwq
jbcnvfcUxvP23Zf7lTEJsUCwci2lzBW+Z/U5pKxmv1bnyFWNEVlOlT3nW/7KQNK52BXnChGnzVlK
qH01j2JAYc4SrHs/pTec/S5PoGU25sBDKi0NdFtx5xuBmx4amavWO1X9owJg8xO6AG5KUsckq5gD
ZFUbuLtxn57YwzOKA6d9q+C7+sjDry2kMs9enGretDFSLEz1f4+w4Whlsby+3Rx1/rQCMNn7/w0T
uizMNb0WFWb46Hryi4sB0BQ2/1EXVGaMW92YjZ0kPvhpNd1YA/gwNJtXuUPBchZQbw9fDema5MoH
HkidugkX9O+5T8rZYBDyqyAYNZ/CVzRmXbY+peNAqWVs05/vlZjQ0QV2Z0GwyYn/r6oqTHu98t/r
MmzYBWx1BI7ZQ2jChbxf/Qwga7TiGdPFnK9/6QVzpKZWDVc8Jn3mNq6RTjMUlGREtK4QeumTmEF3
7rQLOPkZ6WZRvj7S/sUffMoF5fSgvWsF2PwljzWsbXaOTMBY2ZP0GkoxYXzuD7hUu+WcaWg+bbz7
HBqpF/gCGN2XRZ99x0NSWBkgcwGTkf0oRwrS9I6+Xkhu0erScAIvkAQy4itp4nCY1vFQwwqA/hRJ
8UMPkIIdumUwScpyNfKa5cysc8a1IF8SZXW77OZKMCMEIB8/k1P4xFsxrCKAHowD3OFDV4RCHOfA
FP9d6b1u5skhvX08yV2SBJ0VUg6+uQXUiSFIgop8kUaNUToiztaRN7VvwZCdtq1xl3g9Yqi1cw3q
IZueLYxlsw3BkPsbO6w/+PUE6ob+Q36ua+pFh3TP0WRX7jPZuMtft8PGCW49QhRtQ7x0x+1EvFKN
9UvKmuOfCyeU7LiaPaxQMnCIAmGYC/hVKomSEWcDqf78uccffHe15nb8MQFcukXkdewZAB7slgDq
HwoPPuGI9vLZsrVyJSLzzO1iZ5enc9Hg4gSO9Wn0hVAM5DZJAhi0hbJ89MKiy8Bl43LA6DpViIx5
NYCYkLpi0TVm6TvxJF0/zGiAoUOzA6N6JWlMZ5jGEzVxueM9NSUDGHF3ilkAV5s9jIzdw1EMeFMm
+9qLi9a5FM2Kr49GcZNRY4k/IgP50+dXQ5NrLWgK39JmAZx9jATFDr2X783OZX9Yce+CJMSZXuUK
AjzCNQx4oBwyoTgkmIieKZrCRurSEdcyFBXVF5rRhFsAAkL5TufnL6C1mfFwkfK+aJj1q+hTMTy4
tTtANEtWiseYp2z6SVmoFeS8jF2SwfNfkrkysfmD2iP9XUdENnJjH+XvItXKPqFVibuuefqw+IBI
AeMuutsUBexYvHtb6H6bfVLxhM2BbmJf91wwlS+6QIMeQs8EJHMthBVJKFK8mhVAMo7e3PlVrBuO
gqaYBN64vo/NRF+mqsDsYB2JXQ+HJtCjcNXHeKQMyu2TFf4M6WhWA3OPWWVu53oorwK8p7TO/RSY
Tbk0wL0kVm/xQScHyMOB7P8jJhv9HI4F//GmXBVcxqF5CoLLJM6rrZoeu6OuCy/vpwWTZ08/efz9
Y7oQ30dzoccJyg5h8fmfKNFQxIsSREk1oM6mQoGa9B9SdIyskrz084SXHryloxaN9b6bEYYSrTdX
6gRY4es6TdtVulf1sJMB2jTbfDA4tTpABnXH1nxJMVaFVeZJ+r3YFYgxLAQnFMM9BahJcLBUbPME
buRAo6y2vfXHioUXF8wc0K/VbH9WiT+shk8QMfE3wwL17sbjyMswKE0R4PJ/Inc//ZTI0O8qxVdQ
bTLJhq45NaAPGEcqaprdt/SlgInJ127LQTddoM7F5TbOvLgHRtdJlvCCZms7KxSsgyoHv+bPP5Fh
KH4dgvlWPS2oMIeHswbDrC7Xd8bLLZGztmLuFqGvsh4RJjFT7kCVbS1zcuWjhW/rO0SOuRnQdB1C
IJP0tBxqES5uiDcJq0kAhpwb7mB7gfU3MgeCxjoD112hh75ZeUgEmKGoFJXmXYsij6/CKWnQ5b7u
wM2NalL9IIFZYFz4Z/+8H9+4saV/DRyQhpJ0E9A5ImyeBp7IwKkoRKMMxl7+7KU6k7sZP5vBTpkJ
ZIU7wIn7ZjISN3JpVFpc756LvOCMP6o/pdCwouXFC4yPWNXlyfGvoufW6e2j/KYV8dlI8MfxkD7k
cfF3jHdXbCl3nqa13FINdm1omDIAoTlXi5T3kmAyqgGGQeFuZ22By4Olrf0WJM3rX5+bcXDgYofF
clC3YPEdKng6suzgbfkKX+fRtuqtqsWn4cAYjzCay5y98HLEFey6FULBqJ1H7qlyoL89Ob9XXM7N
NJM7FVv5BusEc2MpW0cM/tnXTP5TCUOV8KNv6vxWkhnZ41wCgRPyniED7EWCC8fBX8/qoNZY/8OA
x+FRYhTQgWM8D+UGaG77NxhcV/POk1psE96iQbTtm7iUdlK90Wo6h8PfGGhAgngo2z7JB9XahOZh
mfGhKcgjE+Nvn9vg1JqzSmlO82xHa/MEkWYlaNXNvB5m20pjRnZhUx1CGn/m6kGid04veEgVehcP
7pqTrfCjQKzhr4io1T9qDjscL+kbSaauJNIRV9lP91jNccAvE9nFI4klM/LU41tCinbraHhSk9MW
9oWiC9+rAtmiPk2xkHDHuM7MAOzY+X9iRCRyYeSEJUF7axdMKdjCbWdicbHZZdOts6lKXTQCJdZx
jiwsd5mr83smxEuboOpIx8n3eHyupju/Sjp+v5fetawlC4jtvHOG3NQ2zAMrCiTLAkTB3LuiIuqa
DZ7tDaBUgcW4LjMVeD+vAd47k4g6KZ3JT8uYvoufRZt6PFFoWO6PNxOSzni7I9Q1ZiMkyVqxiVYr
FpB70PCx4sbnLInKz7WKr18+ZRRY/ekUqMXmailj+3TpEcvbjG/dYucdG5F3AOb8+KP4xKv9iHmJ
AGmssgNuFHa3ZzBRSbmI1JjznpMP29+FSRYijj5PdXryk0y/aGZpluYc5p6N7EEdqRoKfHFL6yiV
z/pPfdB2bFUcGOYZ5x4Uix9IdlrXycgdLqwWjpZPi/j18bneoH+vodmTqHo8NKaHnaArOgBqtSSB
wRGEvfF8+QClg72DgPqnXLupe4dkCuTzZgKC0IWWx39tnzqk97eZgm6+KdRkuT6BzVlnlszybWyw
lp/o4rtOtSCswY/83vDvIz9TEJyXXwg8QDSIsucrzgwNZnM0ANE6ny4KENGFAl595P7vtdJC9fU7
aSn/KsOxUgmRryDyzt5AM+8iP+I5HREm7FkQaM1gP1FQm0UyGf1D+Zik0aYvtxwTu3gJmHGGHlfg
0L0LvYPhW3eMvEk1CD5/yk3oynuzFBurr/W/GlcP8+sIo1cOB+pofczm0org7MoVwQmdt6y3P3wW
dDs9tih4simhE6TJJHV6zfsD6f3zuei7WskV7sKxFEO5YhDp/ovbNhAVjl2mKtEiQiMFVWxDcEcH
saEwsOJkfJh68NxjfMFqrGPs8GxKB/cnWLi3gIVGwV/wUNh3mlapHG415TYtGEC88n2cMI2sj0Co
Y2l/Ox1ZkInCUnkICTtPW7CQ6nNWsGGKa/6cFfVwyFpJed/JMxZ9m/WqtQ8dwmKWEWDKpzo31w9c
oIOa4L+at9OifTAaMnHjEK4Fyeo5SH8eExSuPw5F5RJF6BCQTAWXqZem6wFp0Y3RuzfuvbnfZ/eW
6WBw/m5NQbAjwCsj8jJDhR71g8rWe6xxxFulE0Xe4PEgIGij5f8HtuGYa6EVIQccAY7vZuqHnRvz
qT0QQqyzLo3+cRwxWSOnuPui3zhDNznXijPCNEpsacLq2C8GfEcCBDF/9bz6+4/Waon47OxcWcWN
MlZnkihWvlFy7FvUEkpg6YdsmhYl4pDf+C1P1DytUGYHsJqlEWptNdcBrFwAs4md5brH6yehyB8w
cFH2SVOraHri4zaRUwGwjAwiwGQYeswLX1t3lqLYZjwhEFwxFg6Dzl2yRGRilsy5DJYLFC9J+YwM
GWbpjQNHg3KrqKqCC8lqqUsMg0gRFKdjbwy/W+CCc+0ylWumhESdDmRA0oJ4zS+xjQwNQVktMc58
QgJA6pSOCPAnrdsjfAzu01L/Hyg4IuBQVzi8hChZD5NA1ZnqJGM1ej0qmYu84ogxAFn+sUgCC2eJ
aVJrenNCJuu3bwIyhhfZr1qSnwFSvwO4WrUL+/YQsgYVbwspe3mREhNrg1cRxUbvvZav58XnOx7S
Ai/pmHi835qGhPpuh7rn6IIGgHb/ir7tLVKkZ3+VDl6Q2DoRDiqt7If3yNJjzfGMU2AWvx4Sfo/V
WM5W7vd+KpoIo9OBMkZVvXBRI7zDehkME+MrZ9i2qvgueUHDCuVQ2Q5rGZqs0NYBCjW+xs5Y9PJf
VYrY+51o2lao1YPBRB11MkuZeGrEDP8xGMNlijNpuJRsX8XiV6WtJvy9MTlV4fttsGhTotK0muym
z6i5pavL6i+LG278jVrwfpbw/s9MJSmxg2webpFsate6VUGWH43fjuvnukWVtPzlD0MBTCjerjLh
UhUk8lRF9Q6P3y3S9+lb5GyXj1GKk2tpGo8One1h5PSJKwOyQVMIGRjR9YpPLnIAnztsf9Q7zVdJ
N1zm/XyTG5W0lBSt2ocEljTtZwGHylLXiRDJNRVutONc+O17e/+fdt4ak+FjcZsLwB+L36504Vbl
8dx2RfbHeTmu/462e32JxZ+UbdVQrylcSw9nGsl0OBJDCw6ShCEpBHSFD+dDT7rt3y9NV8l0C2E9
x+Y7euiRt9uQyDQvvczmD/na9MK1q53eZEFCcCI0qBRzjEU3Wo64NUTXnBSQyT8yb8bk7QcWK6Fq
zKprToAIqVYfvj1MIzPWfTVkOXQfniXuhOGLqs3FYlA+6Dxjh5rVSoKQ3UUl9/EwV2+ER708Q3FU
9waRgcpYWbiWOk07z/sS1/w75r9bhIzsOolHVXFtrGa+tM4XzPOzdJ/+F96L5qKWIG0D1zVUgL0R
BFqv0rzm4vAUU4Gr4raGsq+wahNI5IDsPtn4xg9oZ7ppoeqpqHDGsu0noLyHEamp3fbNu5EcIwmW
xUXlFOWZ0wigRPuCsHe3OZXtMTXFrcqwD2fT9hZFc1+yZN+IOewDTtJDLMNAPNP7jIfI9j2a8+h0
S4E3UHTC/fLzwE+Ewwd/YWWwzui4tHJbWZx9C8tITqdSgSVwf8qlUAbOXbBDN1Gud3sa3hkr8ysN
aUDFQOOrb60VdfAfPZwpQ0dYlP28OA6Xu0GZA0/sukH674OTCTQtVhY+bnO/RFi57px/pLFC8m3V
l05GnkayQzsvBjav5NfIK0iCKkoyPpN0wDvg6Rzs/KhDUROrFDHf1Y5IQ+boATRH+cLynxz/VJji
e9w43YmaaiDNiKVJlzxW9HUlzyNPrfGtoVPW5PKrRKj8NJ4Lak2/zi8NmWugdvEt1fXUzutUhbnB
6oXqBQDEKo2FDEcF+9C0r9NnyXf2BTSZ9q6wTUvEv7nUCXwIzET0PrUsRVsbe+JbfF6Xl+lER2+x
w6Vta61IC3+tUAaUm4QPHwDk2MBLosVl8buRV77IWwsbG/gOp4q7L5ur021lTnlPs+RlbpAwLEF9
1T2SImXWzEWGDdt3C86LXgAfW8uJy5YD6ZPWrtkQdeN1YH2t0vXeObrFrjXrVjDM7CXD3g1StmYT
7d6WVkomBGE2a+wuoZyO48J6bX6Sii9G3pABaSRP8re3xdn63RgN05LZ0TRbUoZamaS85bHrOEKF
2NrOS9LYD/9fgVN6CCG9BbuyitrikyJ4sjP1wYWIfb0RqYKSANJaS2w+fw5WxJoTW/yRzXrmX4pL
Tmz6emDaeC8Khgw5aN9G+uENX25T3iIWPI38raMXtSjVR68xNkTgfL/4G+xludP3Ii1UBOhokVS/
62uw0HYyBGF5WC8GdqAjV0KG7oreWrccoqLn1z3L7MQT2l79MkW5DTfMiKERNZJ10F1UYR9fVQJq
DGD9c0+jp5ACGLnGrnHKXawlS2/RgKgJtSHLdC62RAIqlKzdDzIeQI8EoCOIjWcOJk72fZiG+oXd
dd/3JCttCZFYSo3gDwc6a81OCDm1Yf7Qs4NEgLlPg6mL9JpNnWEMq9iUMZGB+VMSxgEA1j5CUMLY
Foef6G7g/PZs3vKkIDXuBlip1m/4c3DoalO46GO56lNCvkZLpjPtO2j/rsXe9rBbrSw3oBn3CouW
8ro2UmHrrGUtfODT/HsNSeJiwMXO0UiPxVDscrpkJrlG4oP+pGHd4BgE85MRqtYMn4fI52fe1GQw
NW7aJkASmiePTho48aLxghiW/h2EiQkNLs0Tog1YMTYecpVCQ5ZtfPDfLXSVsq1MSKm5eV4rK7EK
GJ+srxhx9unq5YcMPq0K5NwcoLdrsazVYXuNqlIlwIoWVVuDL8shStcDI9R6DTzfYJAgwqt05Wpt
WF0F22moQ7DjtLepKdYPKyVG1sc8E1od7RG6/3U+xaqxb7gEbI9Te2BzBYU4CzME2IiEOUtsQ49x
+iRCHgOuaKJOfBH1JCm8Tlq9zL3SjBzRdV8zEWHSMYfYn6MoTfra9/QkAzurmxCPmyC84E0/Xa9f
4Zjt2hDPtVZ4i9qUNBh0WXEyF2eMzkgQYTLwOk87AvKgq6QAKwyGZLPTDsdRRNvi7RBIgK18AcUC
ElxybugGeRc6wd6Pt+rAmiUjCoF0qg0jDKJt0eOhv946S7Eb04QVNE+lAd+dSzVUZmqR+jRviu+f
/0TOU+nHv2MKfkTLIjP/1J0JSMPI+h1tQhmtyzCCaxcisVUURaCSTr5xBb7pFIRvEN9GmlHKcNrL
sRDYGwUSRhPBTDGoW7jX3/QrKTre+ppuGF/LpjhTLcqFeVU/f64HTnQOIrhhgwWKgvD1kME4V31S
6iP8pjvQKPsstL/a4P/EscHOdfXWX/55brYq/q1laDkAq7qfGYFnJ7Y65LPt/jjKpVo5HZOvISPR
qA9eLAOgXLCuqA+6V++YKo3L3JxRPZ+jY7joUNVJhUpBQowDX+t6vpBbVQIoR/vU6n1HEoKwIUzj
9WsHlcg3v6DwjpiEWEXoxsOBAmhC52gVrsQrTCgo/CV6UmqeVzNBLAJyJ2OU9QC5KP4ziVimZCSd
6Be99NC0GoJqYMslqIYLcwijrHvwar0/xdJytYdPYmtHLxSPDJofsagx2HXkxTaduggW3haZsSmx
ELkQ8SswpLzt9JSilc3Wm9gkbj2xj7JSUcCvdy4hs0fAJ3j+9GcdsHglAYxjafMHFaXBNlrJsxUX
ooDrIjn1Pub7PO+9DI5zrx4w0vUDPYAJhmHpQ5oj4plYR5R0Z5dLGMHyZK9JsvYwXmCdAFk41xah
gSgQ+zx7QeeJnShO3FiH4AdjHYHStyd2+UBSf1GuqCnAMt6nS21UEUxw4+HHE4OZGWbkx7kpOu6C
kvob7odX/QCBDa0VmOdkpTYAFggK7LbPbQyxkE0pXWhfI9tAZEhW7Rv4ok3Vi/dOXCRV3YWcd35n
/Ov2Lh93XJ+3SlrHc0j9/oZBoEtHDnYzqg3JqnPvbzF1+xABFWqfitCs2KV4S9Jg4Vr6k03JPxq+
3bh0Cq2FNH63dnySh/rD6UAfy3DCtBc4ciOyS4Cr8KbsrWMaB/f2IkReASY9lIu652OiVRwIxHwp
QjYPJo5/qJU8X0sdz4vty96yFIH0Czp+/Y+xwwGzNMz9Cao47JeH1MMvp3w/bj6/HQF1lO85ScB8
EKbL5bIw90pkmK5RDaa63EbBbuXgx85iJxb5LJKrxFGzj/n23GdpA7OAdTnFHlk2QXfwyrCcl81c
Lf0zgv0Li2Wmjm26CUkPmdSi9KQAYz4rwZS4r984zI8HYWtO+KLDwH3C/Jaraf9TjVt2MltQNSfU
l0omoRmOoh5tMQ6u8QckXyn0RVRhpZwGS8cgiq6JE2zpY+grnL/FIXEENV+aFj+DggjYMkWCJEdR
eTUwMvEB/c1O1G8NZ0KbF3nQTTEmh0YKhgTpxv8GJLaDLImfGAi9alpGheasnU+jFjog3Q2asJVd
meweOWLscoSnesWpHz+Ol0pWOQrkSphN9ah/KGe7tJL1Hv8KJ/s7bPMmyD96/gJwjEdcn6RVZM0I
jwafcom9/WdCMOfnaK8yYbW8ByGi9C2rqzVJ8gW935qIEWYsX3Fz+7MId0kmFwJ9zqhIHVpiOUnn
Ct4p3lYsE5qIehts/+g9craUabgE1SEhKOwR4xxOzlnxGAWP4bs/ms+C45zfn1AadQrVK6pr7Lhw
sRRjvWh0pcYDDXkwcJAH2DSuH8esra5l59M/N+fFfJe7CC7DktELC81T6q3XhEjIdLU8ZiMyjNvj
SPONMggXbvNUJ1YXXVvcK1l0chHZSoZs6Q143rEzOPvGyjuzTjmiEd/7fnQyZCvvPflSDGXvZsDF
XgSFiPCS7xAS+ZpYd3P8MGLCHwZft8E3iVFf5lBzP2Dyi1Piiy5XZwvdH0Le0jtLpM6bTYQmz9ku
0acz19k4G777HzmGXbwqtrk1O9FPaz4UpnaJZjsEtlK+bCtzB3cXMreUvhB1eyJmF7lzScQ3wgjZ
801I0IKbeJoFS3DrhzAwIeh/OV9oMYY8hlNUEF0KwaAsNTmUjfJkcQQShFy2yUWeXSgObufaucbI
8cwttvrNcJKPikl4k8cQU2lIQZ16z8LfHGRx8i0omny6/mKpEEBtrVaswWl5WQUfxKdUrIUe6XWl
ocH2Go47RvyBrkOl+gBJQc4rAGf+patnUaPvZ5zHGP/y68xKvZxCf+NW4jkedp4/rnpdWJo/IHbL
mE80zM1iBv14lKJU1OhT6VzVdLduA+vgHlFj2kujrSuqFYuY2LDT5F6w8Fb1ENXz9WCP+h8HaUZZ
kQxabAZ2QaKJl583ACqvUNDE0hBBI7qQviBOLSrRox4TNwW78ZMlVhyMVdDK4m3N9VMOKSaUcydw
yWQiAtnn4ZeP5gIBbYOtTsr+vLccTtWaH0jRi4Z1V2GNBTdpz16mO6KESX6OJzwhVAAKYMPL8qM7
JAV8IZmo3QQbaJtNe11UTzJcdHOgSEXwxZBXjd+1MSFL9aXOeDlj6Af4rFALAzzMS4qh9HJAoaNJ
M5J7/1aNSDF4f3OJguVqwQOt8+solJg8/bcm93vD1OMQdYOZNcoTsL5QdBo2Wg0mEUJ3p+dPpztT
oBUpo9dH1yCAnpXXuDv/9yKH4eT0KSh6jUBeoXu32eTNxL+UmrLjiEC6uMlorRza3reJlHFShgwD
NJJ/yuOq10/od9dXzIUSpc6u7E/o6/l7YE3ra3dAlqm/k8bBI/AcjvpAIyORF2guVlYrpalm1OvE
481CmsZWBzFCNHDIgeG9YB3HsLLzrFJGo2b0OL6UQivPnLgrWvc/1MAM6s2leDJ0vliH+aTk9FRF
pSriaBkgIMJwQBS2TeHT7XdlQBPQFL+a7J5v33h6UoL7R+UuvemxriDd0T/IU/gOXuzIKmImh46l
DaJQAk8wXdWBIvPG8a2eup5T+dKKwfx+hEVawhzInda7XLNLmDdzxYzkmtTGgliagFgzfYyfFqNA
Imq2og7mckJ5hBqSRWXtDqMldT+i9Is3WiUuxFRPcZr4sg1sA6ZimC5Q4T1hh3YuzKYMu8yVIK+G
t4ipq7v5tfply1kQIwwh//oBpjDfOIvaom/Q5/BSNKKptIw9oYY4nnSjfsefI1HB5x6nlhfWbBOv
EU6EeAYYsGDob9S7XnGi4rB9nyxcNe6EbljjRFAUjnPUhM5Nq4N/v7LcK++uwUc+f/rYnfZUYmH6
x6261htzt6hwoiMUovIUP7MOIloOft2dxPQFJnEuIZReTdIiISZR4NgoN/5kw5ORaSlZ6jpTC6At
UF4gMC9nXfdAgBxWL1xnuQFUUYUdWZL5kiKVwuqIlTWmIlkvjQiT86FWH9WJDIsIQuSqens6P37l
RAhgXmfnGeuuHaBThdoWYraWbMcq7vhipIY2+D8FEVfCbIgfK4970vSk5i9VYNP+8WahrZPEBEhx
kqu82QuGkR/08a5JdSpA3FdXSiwtQVnxGpjRsUTnyingRolbP91USvyFMH0oPjZVwltviLud871J
rPJnPClZAKRvLRxy4Ty8lP0AmNn56h+7xy4L7RqgjK3KhTm/MmW9o86tc67D5UMTCbPCgT5YcKGi
cahYe68LacO70siDUeTgnD0/DKycQpdUNWtw5TermBTit9mEbLRKKtP3s4d0VTqzKiCic13HcjXU
pLU8SSDqAZFj6E29cI2oKbueRGhPFZzJAQ+JpXHAzcuf5P801ibZPDuFpLCLsAyUXyNChwa+kz4f
3BCpAuUUG+1QUF4f0Dj4B94UmzKkez2TnX2Md7cGmQxkA1eSaB53E52234I4pl3bC8ORWmG5Nyg/
+8TSDSlze2BXH6arK4ScYgUTl4fRWmc51i8aD7CuUCEG/98cvaCw/33lc0vDhX3XdxXKPlpO8bqL
NuSq2vae611yd+YDLCUThTApQhQ3HVesOzO7ugR6RQrNrqoBToB8KwvMyRwdvCRa8SGNCzLsBxmH
NByJEVuuwnEQd0mk0YpmMaFAprMHcE0BV2TqX7ojF30yr2JmXzkqawvXuQiMaGjB8JMHMAVPpUTT
58GZ+I1b0gsN1YKp1M6uOe37Vn7fUV57ses1NzHEHuKSG8MdyxDa3ruecjqYZUQw6ltqbB5WXeUP
QTD9fHO0KUUkg/UV9IoK07796MUBSTxbdiMKllWpk20liu/D2KDDlwrumdftu4W8SwJPznnf1igU
apSFy4GxYfjIaAYy/QACFHFxegNnHjaHw/slAn9L8fksrB106UGqmrfk9XiAAxs41uXytMidoLcs
4NLIHiRg3AHJhwyxcrrxpFrMNrnJrepqn7jOCU2MorQQTsmHdQjadm6/1wvF2Uy5lZltaivzGOyZ
xnF9nlupZhD1zUcaYrTjbdMzlJUYyd1cndAtCnFKvGtoPmCtYmSnhFF0c+buS3rYWsCUZ5CB+5c1
kJnXIbLHqmrUR48Ams5jDAswn/L1CsdP6EOQL7xizcrgsao7+pQi5jEd/PG3VDgWi4hcArKAXi+w
nPI0wBszMB6sIn9Yn688emB9BC1J8xKWyqzxaG2t1j52HljXWapUkT9uC9EdX7BSu+DFLYIfsfqP
eCdOhdfI9XaBizjD7TeFKwg1vV+wNhuKePlvFO73AyFdv8e1Urqh3BqFUXz4eo//CD54oYswTFgB
HXl/Jv9gA/k5LW+Qv/GkrC+18ajv4rJYAFLoB0FojA2w6bpgNVivrsntrOGjZaBUYQ3UDBa6p4GC
6uuXX/f55fsaEEJG1zOKq6L55dbVYdyZq0aYlbQ7RueKFjuxnZcNJKdsaD3yRPLmqMji/rjxbfsh
vczW2TIgrqIBgGtYrIr27DVcPV8ILkfj/J3pTDzjUw5XzzVGzl1hh4BGYSN7W5u5VepYTeCAISNJ
Yj25lw2BxAOOkTyVxFaQkEAKTgIj0js+x2h1LHUrdFVwWFRJBv959gaGWSW8Kznqb7sr2tYZ1lFV
FBOH15SFtmifxfj6JvMQAzj0cyq5INHwdh2xPg7CSWB4ikYo1FH8tGnPbGFjx1F2qUmJ6vxjESOO
qIFdBzSU2k/EdNCQnBiNuJIlyBzeOtuZEkbsF3NSD7WaubCUW6Wb6TJpa1NBxz+Y17Kv2XsiqVZ8
v8nwly0OecEqOSHy0H0bgXXWTVZ9EAwf7ypXit19jnXzUMEaI7O8cegSqmYLHgCT1RWU7lIXRSTW
yezFO/tgCyxltIqchGd5K1I6wSpzcdBUsK2wSepqcDS/drD9WMER+BOzCL8IbIicJM4I/RQXzBUV
IOQpigXl890qhcBezKtfFmASbeQvppmCL/981NuJDcJNED+XLN11A0XIokjiVkOcYBmCY6HMrWhT
l+muGKym9qTKHvL7cGGxq1hshGGSNmZ69wSWPhsSTHFd1BilxzV/BaDMbAFg4qpAu6oIrZrpxHVE
eyZdfDV/t3Kvbgfl4RsZMjpvcNTojZA28jjiD0myCYdHSDW+t3jdxSk/OB5ClcNwyrpMyMpXGRgq
lx/UwBT7Vwm2CYqdeZOh8d2kdD/8sXj/cKhH8pqzDyVcwqUj9jGFs729uUUvlLY7fih5p1WE3t0T
AGCDeb/jrLIPCNRWr/ZBgC9ZrfCDdlyO9ylQjHKv01xrN8eFP80QFNQDRXGbyHa2TiYDIkSGRjxG
7auNIqpRfE0pqHQFb1l1ADZxYQWeJlkyIg390JNpl8bDaXYDEDjQ16LtT4KaTzYViARpBxj1RpWG
ZeJHQnF5MT5YJEXv+GE+giKEn2jn/ezRp/fQ+91Jyp2Fl+GkLotrOJuF37xg8KbGLMh2Jhrx4QRY
FXwydf+j/UkCxS+kgrbOccg1x8tBOpPli/PvGFToURifwpIQOjm1A8WTw1gGjrVckry6PL/eV7Y/
s1PdEHxOkat6Kahfs6ck67CMxC/cZYkGEKCQ5lvEvI0QhXp9/DgHos7WEJtmeSa3VTs6Nv/jJPXR
63YBrmaiYAzYiXBkE5Dr93v5f76Dhjzh2ui6svYcV2oBiUNJbQ1z0TXbpxIdNqHgVuW45FY62khW
hLP8ZKcuP1jayZ1eR1eaZa9yeDcqUHfuzH1uoX1HloC30RLvuRF7rKU6w1pkbLgeERGiMpgtpcyl
HxNiV3W0I1ME/XMWviA++JU/mky8UTUuU3RFqnNpGVAteIRA+tw4w3LCUulbVegfxS1agb77q51G
oQTYz6P2EeJg7/aFKxXzBdU2X5AMUssvZ+xv5TVe7m14cY/GmNYCXZTcqv0uOlC2AQTkLttmuGgk
boQRPmIAq2fgE6zAsjXsRk1k6Ek9YRNcatIbaLvuNkoEBnIOrzO2XcH3eggYSlpq7lYVZ6A5teor
Eu7ahnODPZ/dskBxRuR0j5dBb3kJhRrHWyzIaCi2ouMO47vygWSdx8gGVxw73POdj/sz7In5Uxyd
7yvk5A75Sl1V7Uils8wb1Ex/nDvuUhbIYu/nGmozIUNHqk/vCHH85UygTtyuD1I6N8FM4ybfwJFn
ZGSvLBAiI/g9ZX0opKCnR/bxCOBw2hXqLN1HyC9MBEa53CXQS8urMP3FLw46hq9WvqBZrJIaePDh
TWFGq9smhkJXbR8oUX+5qgIZyCQcm0Ilxp4gDTQXWGJCe6Gkie8TJ/XRd3BVXxMrJzk8kbibe6eY
D+oxr8gGnw5Qiv9QcBxiJ5/F1tpesAHxUzB0wWJ6832e/E1nhTnBLi+nzQE1WHnLg+MoXv2zqFoe
/hEr5drrzMF+EDNqEEiv0zxs5Hzd0bqOt4Mdr9eUlK1TEgpRVpvPcYNiqGLMaa7wzNNgJKmybVyR
u6l2TGGWX7KWkBkNvXGEj8oEzBB1YciuPglyj2jDPPZCUmja5hOFf+DpU0Qydli2hSjtXrdgBTe8
hpCAhhVTPK/CoymXXMQm8Lzo6fi/IFi+MHAuO0BLxauW7PkhEmKHqLRYNo9mFoMX+zgZLfXrfzd3
EyCp+CphYpZKjJNg8wnVeOO/Eavtj3mdE7dXBUVCY/2dQ15Uv7ENxSivdoE4ylQbCJ4ZxiMvggif
VaZJXaje2aBfYXkjgPZMT2me7dpeK/FRXW37rxjWuiSvZxe3iy8S/DYTSdYJr1G63DF06eDpiUeq
exf+jtFVVASswXoF0kyvOUYKdtQ9RMJviqhLKFAgcfPMokNxMTdO8o/XSKadxAj+8Wv6YMmQol6F
kQ3pLqFmbxrz1sl56ZToZB9rlLdurzYCAO3EvtRzQJQ7FSEVi6zLHSzgHTfy3tWD8r7dF3PgS96q
cHMHugZBFruyEtnsehjIyKt/kdIFhuAClYNrAh4kRbiLjqV+VMQzA85jaaenfgAs2LwBxHyPy7+j
mlB4Pfy5OMj4oSOB/3g9hSl2w49B4mYe6H8bkyAHWntxLVFA7+9LprU4K7VcwXKWMEjHM+xoHFEp
RfHkywQ35zkbuEBAD5m7Uyv4NZvRKy5sYIB54Z3wnxJDupqt8FvU/iGptVe2DJZ62Zpb+ErQWwmu
r5/QQRrr202thOu21d+k4O/UeJbnYLuaaIoO68oQnA5IpgwV+qgYGmf11Q5IdaBuN91fU6mTlJlu
vHi0HJTjudjclxovhTqNcKAIZ5jYInqO2YO1fimGcWykkna1otXsSxJY/2ayE1KpsHDz2YQykB5W
oE22xNIcbevrFumT+ZvBKWGgWLZN3+isNR9GJP1nM8TRec8kjAww5ylwqjI1qcdX3ANtPO+bfA0Z
8gfjiDeZG8cWomQJ+BNgT0dZbDIKWE2CP0mxbeQQh0vFxrxkvQfviKF6cOyCAw6pB72diEa+089x
PnlwR0zDoe/UbPVB/fGMpEIaYxacYOCdkI9RtWOQJmQTVWu5Hf1nZqNS7xlTbcRkrZtWKF+hx6e/
ch/dBmxOb5sX7tU+rRQaYRXPn2P+t2cMC3rkM3jCDz1acBxJRffFTUqsNUaveVKGLXsKmeggSgGd
KzVheLZ70UE2jf5OaLLjrgxoMkrEALTIHyeS9FVlLyvbuAoPdd0fgK/8C6YjVc/tjv240P6mo4kI
A4HwLqKJB/sF1aMcERDxeKnkwycFwgF1EB8mck4Rv+kbW5OUs6/GGDyFxWYlnNIwNZIMHQVFa+q8
3FIfOgM6qOtfoWKhqESDGA5FsBdeS/0BEDU3vqrioXvbIwOaTZX9xfg16ZwYSa0sruNLQlJxfq0b
riCjdljni2WIReMeqmLZmYJtPKgcanzjXBCwXkAfUH9LPIJunVN8a3EN6GwIpcFZ2uJ5TGrEr4A8
n3LaA5zxEVj47rqCkyWaEZsV9Lruf4S+4g/mmUqSQw5RMDydwbSIRV40VH5+emVFwt2CmLMWfzC/
vdYaXoEyVAJe2raLUCm4+97GNyGioAdEI6+ywlmjybh1qEdpKe+NmKyrDPk2b8RUhZ5MkWyQvWbi
xBihcTY3D4DLCPFR8E3Nfh1OkZ5hmHdCPiRRhpnUhIx8TMP9MMEsOY9khdYwBQtdCKA6nN+NGOO0
ZdpF33dALRYnXBBwJ++f+iRw3abBQ6XXaCw3tIAc0dNvfJ1O2SU06iCkHH7ZxJMUQlVA53Ksik0J
6ZR/5GlXtu7Ewb8T3EOGAxt7xLWCvG/XjYEf8OgnNEFUXfFK6WtyNaYFJWXBbrvJw8ieb5GmVn5v
juu7wSkZSpyCpMzmEEHY58QRCRcXPqqr81Oq137eiJXPbiV2B04Ss1EfHcfUuYAk7hHRMZ9vYK3+
JfP9VJlY/Wrr0KMeR4eje1ETp4PFOEnCoo1rFsTpEfJ+u4KF1TP1MKDwcZ/UWcwXe1ILERxAavlm
m4pqAi/yPYzg1wjU6uRn0o4QTY8RHUUh64lhRLPJnNZhiJTlpEhIh9kC/0Uc8eoOM/hktE2Z3fZj
VFn8o3ltBZy6qbb5VpHHVKFrcgsadxKI0UF4mIsCFiMdBgqbM5kUdnYDEYQ87MmI4v7eeo95kBNJ
oSGYU1PFjdBWOOuYKJrW+wh3A8t0o+JKk50stfwnbUL8DwyUxwQiko+NTPeYaFVaPHvlsTgtsLBZ
vSb4nLT0tVLsfL95/J8oV7n7FTZqA+ZVlbwtcVgMIWXNne7M82UGJFjG1G7SiLrzyddC8lh1GyM+
dJuxX8Nlr6Si6u0dAy/edIDMS4lMdcYgjQRck+v2cVAR6b8mFPXwYH0REa/AZMpg7XjyT76e4pHw
RWiz2pGAWEg654+RZCFMBqugDzH6Ge72qhjmRssRBaOdLrLH6TFj0qNsVfYKXAbFvFWnt4EbYMvH
VkZB5MzAADxsMG0VjkCTumQxdf55TKTJGfg5vdL5nK5b3PIbCBuqS4l8KiPd31gh/mtHrzvznda1
Qg9JpzlADD5Cb+71wv1j3duk0n3ndGti7RSQaQ7Feh2rAiCm7EJNYNwWY5Uu+oZAF578RLPztaLM
X9hbeb+STSkjoLv64UpKtAXhqhaBviY8jmyfY9mM9TGxPitJDncCbplwjGCdbiG30uwtCVzNaRPF
XBBP+NYqyMT5YILflfoRbf6fkVMbBS6maX+RurWfCjgm7roGEmVWp7HQIDBK+JuCyTmYxm80lNrH
/Ep2ruTLb7VAkRG+kv8rz/c8u4Qf4VGmvRatvdzZbaf+IxMI51Qh7zoGSohZNDnHVI2XccsAw0iY
0vkT/1JaJH9MaQ8gJG8mSrpcp7ISIYrohxyIZH6RHVJ+/12PYE+gfDCMpM+q+mw7qyhp0ufuvSFU
y/mUd+kU6l3mh1ktU702UXpOmq6NBCfsiv97SJiAIfmecKHP9tAa/IGy1pHT/tcohFsTbJ4xfx1A
mE20QcuWc/Vfn8hS9QRAwOtQoyPHcrj9k6f8wr1hfkb0ndpwbuuBD0TDkxVrxCkLkSUJieiS19TI
2cu1OKFGcUcZ8CPYG4AOGwoGiHzX3RqmSPRrm/xV97tVMJiRfD+XTdReMwYf8pCR7GslEXLLnMjO
dHHfqzEv/FQbOj1E7MxsTBoe3lRiNqSDT7Es0QvCW/Lo3/swXLHBAYcg6BecoWBXmtZCIQQT+n4O
sg41gSIN0H9F9NbGryURBt2sDWjXnNQ7vcV44Hde7Bilb1mMs0xDY6abmvl3p7LeMoyCrJwN27g+
t/9gfac7VM8MgHEi6X7n5yR2VL1suxL3F50Wo2YOUstmpJKorA06m+DjXDGctIdr+rAAg1sNJ3Fz
rsTGnfIKcjHkvZ67a8/KMlay47UUXPz1q9GFxtXc1vI23lZvldBfgjwAHqn5q3aRW/Vl+IT9cTOV
elpaVBWJ5WTDxEoqnloNdpC1WDs8KrW+r4eI4K9wrKSNgAgPCYbKfMaNK/IG1H9ggOxx+aqt14gu
MitpOWJYNeWwoXWXjbzMzND1IpEjOmx2nS5a5akWZ7EKgo1qum5RdfLw6v+DtBNAzneYm0x+8GTR
H3f9rIn0XWGmLuhdG/3ML8A/XlXnS82Dovc7mck3AwlgIM8hmZtXIPfYlL2e0C2Ce+OMrml1fqAl
L6AVCdLrxj/uc8iuJSWJrZs52At8EKjbSShEWnZQ984afsE0DBcnrK2dqU4ZL00DD9qHRHPUYbsU
rOnibdu26uxt6zEZX7cnDZe7dRMiPiqr3Wiri5jkQsm96CZ7xj7Bh+sAnePwZIsL3SIJYK9K3HZr
g+1v9M7K4bL39QmUi0iPZ3y9CSU1yAUlNKhF0VFWAHJQEoA2YhkiPdp4NAid9KiGwQWcjniH/5Fy
XPcplvH8mG2FKYx4p++q0uL8ONa4Idvikxv9JXQ4TDrDi6IMbq6/x3xfaoUaFcLl/WO3pVCzW0u4
4zbktyBMqdSXjSF7VGKN3zIi3FZuMMYvjmnN7LlfV20MxgnFwh1ymratB+PjlyRRcGaJxmZPh163
wVQdNLI/hc0F/ZHWiuGeM0lMdsz+ff83UwKmdVdrake7q0OYaNS/DqBB7/xAjAns+7g+xMWV+zSN
FoMdHJtb55vFJL+kbOEFZJAW2mQeqEzYS8VLRqtvDlCTq5610j+TDG5ZABP5eViTsnBZlJJMBxv6
uixJlSViqu27tNAhrxVUXXrzt7VeaxMxrp883CqKPA86+ps1+uCf1ZOMA4ub0Tw91GJl3ukQEC0D
dIgDc4kTpx459IVDqoorKGUSBrb9JsdusuWIBME08UvoyPzUnhucZaKQCmfLn+AEJTT+5RhM5cDi
xHycumHfFxa4mdJ5zAolsQvYLWKXHHMlFFXAa4xHk979JhKOLaLrUVZi5cJllSK63jzkBH9RpVAx
O1t7uLGhiJl6XN0WR0CgrjKLev62EagJd4+yYpVz+JUgsGPgfSJJZpMPyZoCVVoe2+MFLJyf+AN0
8EHo51+9fzxvv08AVbaAoJ7vZAE3AXKh7+J1lJs8w+AgQEjJAIyDSb3Bex8UMCZsqC7j4dXjiVZD
kaBn/fljuUm2uwzIEy4IzxHgaZXE3mjwBCoDfIX3fWK0Sheo9GVJ4nD0usgIyWCPZ5gK32Ei5nFI
YNsX9O7cBHGorPP7GXZQKCbZTO41yet/nCbAZUztJYK0JvGRmFS5CpvkjTnOp+8KCiEzRVunr7Wh
EfDnMkFDFtFwub9ffNmKWr7qm+Hm+jFKrjppGmPaNYdFuNb1zcCVzqbcOfkui6pVOxqpbRwf7hM3
gmx+K9Kjs9+q1BAq63ZeRkM/hrsTJMlR40aHpduzf68/YKubb6vfrNTRmPi9Y3WdhtmNEKUwa2m0
YtS9gNyIgaJVD3RdzsjgsEFx/kqsfvIfQOCMe5qRLehEuCI7DRC4oyc4I0cTn3t9LdWJt9SCzc8e
K7ZGbfPKuMSYNXeWpafK8LaEfdtjmOORzYb86AzTDOiwngzy2kYwGFtbaW3DTX1vh5N74B3enOn/
p0j3mD8bOr223IkIFKiNzZOCXVxp+rq0/W7ikR9u1esR0pD428KqhyxXbhlrk4wt0Pazys94sFER
WKW0Pho6Yy0e3WMo+VT71UWvnLsnE5XiEv1FjPqCaHnhFJHsgrdwElt/ml1IYnI/amfo6AF7LB76
ZJGDfd4KzDokk5mFl7nEz+PkFoHGvzeQSOH8zYZo6lGE6LH2FtfXLp+5iOm09/ZRMv6NDhCLYsd/
bKw0mL87t947OHtOkFRynmeaKYEMxe1LjKOBqromGg+4zS76hntnREiT9CPqc667jJ78XeSVQ0X9
F7WiH8a5ERRekfMZjjGV8QL8FWwoL/dDnoe21Q/GDQ/AqbI/3JrMtiapBtNaz37cdCX1ny6iXtUl
bu/dcp3bCUfdM5ic40F6ZYRRl6COwU1numsH7qyW8HVrmA7ewdU9jb39jF9cL7dv75o/17d0d3mk
h0LvXv8nk6M084q3vU7nUUvQFcVrj28/8H598u6AFshGoCV/FvGT4tJ6t7NOGkYG5R8SyQp5zQSJ
GwyJoJkH7NfwF36hjqEuvdI2Dt8B2XPfotJHeiRgJ9igLhaVZlJLNtSp/zk0EqGk3bAkbsSmqxG5
6lMxgerkTfFjc15weLx30v6RZOjyeKlePnW3DYsts59sGZB6E+62iioMdcZYCfHP6qSMHqNHAgus
vckY99/DlN+DLJQJLPIWSd7qFQRQUT5HPf2+AOfi4TV4nxlL8GWte+HMLcgrv8mYF2OWDJuXUdsU
aK+jtkJsqfIw6wmXAbB7XKxa9vfCZAgwCd/yGTJJKhUX++z5fhTYdIrbZTUPCOVAJqB5NqmNmJZG
oueW43lc+UDsg/oQLdWRefslB/H/Jp4SNXAdBmuLPqL5mQ2qYrZo/i2qmfHClE/wr8hzXN5y7mua
3PeryPhMTFaQXxC9Iec4VFUK5oVBP0IWBHq15zMy10LgCE1ENJN0mDGQjN9yRNaJgvQ08vb0J6pS
K5sS0fw4fqGIBBC3skD2JXJgwpZdV5KDG298GgdpsT3cfwwbcXzHdhJAjQdK7XKBG6FlJ8olI7xR
dsupv8xZYvSMZk0S5ECxDxADp3NGPvE91twuCQWZ+WssIVB9b57U/UbO+cS2S8uNVgBCi4Kl59U4
3p7A9XMGeKfM/vRrMIk7JGDB6HoCJJsu9ZAiRbtbOdy1zV3iL4KGSLIWw6SRJRDIBo5nWgvs9x//
spShRngu5B/397vVcEQJdRiWClzfRFuuOC6vKuY0g2FhyVH6GShmtNt8WwP65k/ltejBZwfUOqlv
Mf/Q0j5f6tU/NHdk51mVgv1jTVqTIqBpg2q5DmAeZJbco4laKfpL2b3vnBa0iH1I1ZIf5L6d7eAj
gSL4d775rTQ10Fh4VCsTrkrgotcWbRjdaCasWIluKDsujzPiT44FP46xAinXH8ZufGbu7a9ba5i9
KZjhRMSiWqHPr7mu9DUiweuPWuFUOqiC7VMddiAgW90UHsjvnEM3GYTQMWQwlYHKIaBpKJLrz5El
dnN/Y6tQ9HrfDWryK3TM9aoIjYJOPY5NZdUaLQxw0iUiKCEhzT7KzG1WKfmBe0LwqIkDvLmiLW0w
oXBwfH9Ri0/H5JKavATZNRxOT/JKap+xkTozF5FieMPmj3ySuCoYGAfrzPEJ7GG1Q9LqaUelqnWL
icO7OskT8IMtg1U+VcECDgU5Ut8pHq5ECCCvN7VNegJlDEcEX/VU0vTNCY4g+RuyWUSF9uC0Vxfb
mvCjwuQnWWbaTSiqeZGMJxELka1e2ytnyt0fkuFDNrBz3z0UiXBHMwNdKY+rQMSd+KqHbx4DZWQE
o+/HYQJE4wYW4claMWMUf72qMEWUNwaKDbQm93A710x1v1pX8ucj+5zM0HInqrRBv/AkwymJ74zy
CQ6KWcUPDUaYXG2eXgSlmzOrbTjq5BXb1NzLWQ0/5fW9yse9prkp1T/KZILMbEKfqkLTCeIwaTXx
hyTYZRLUe33gRik+8UUqZtYTN67bSEYLjAElhy9m7gBs4f/3IctC/hYijtJjP7bEzVquYAnegOLo
clyrd1tpoIFe/XNBXde9lVqCjOcMEiCWZmHDHtlR6om32RouhL/UOJfzlaL5lFegkwWKyHeioVpH
wV/rj4z0zQMEnkdyBaOWQUnDja7o66y4hDo6yyFy8yPW6Rbyz4v3/2uH06C0A2C19GnKX8u8yo+A
MdQW6115lfJpIDUKh8+l3scyeKjErPx0kmXITLMkAXp5gHFLxIiLfEa8rKGVkc4P8ee0HW7NY2F8
DVdbXj+DeBSIEcyzXElqI7wJB6nQiiUTkFu3/gzDkAxemrp0qvPKKl2uWMqDtUypqOfxKaqCRzDK
oxb5FZSZikAZy1GX9ioGefHbOHKs/oaOtgG0tNG6n5T8neFjy+cb1O3BSheQvrKBOHYrf7Bm7FXy
DEcdVzslpvNb9A9s1pzf+7uuGMI024NvcvJJxRF6qab8SlrT0AKC/qH0H0lztGsFVjlVOLdoEVra
zaezZY4LCRWa6QSDzYxI+H9UMRIOLzw0qgFz8DO0MTIAUZkSk0gN29e+yfSIWNZUDeZy2NqQKoaS
lpRNV7xgX725ZTIwNOk1wubHllM1q/zVqYgzo2o5eVNK8XuyWtPyNTiQY5VwQqtL3rV6uemzCne6
Akrgaa1oEdN/16astDLVUrtf748cxX7XHJbWqOI6PlqCYkTd85Ht1dYaNcNKO7oTdt9KibeS/kz3
kdXi6n+EwbKFQRVPys+b8CiJjoWuhJQXOf+dSPNYdOninyAHJ3DSF8FD//R2ZViFdMqRKVbmgzYT
SON1XUoClIMiYaczIKvaaUMeRgLrGRZDL9U1h+QwXWjRVX5ymbLvdQ4zWA3yf71+4NwcRK5TGyVg
RYD8gzRqSjv9aAlWA54KZ12y64kP2oqjLGabUSZ/r0TyPm5jfOm5QzY8CUIU53lyIIoozQbhtUjE
14ky39KIE+638geNCSDTymyLibe1odepPLwO7Sx3ZNoDlzgf3hrM0A0Z20J7t3U5ysTgEph1Y8Mh
3EfjD+lp4plwOwcl07OXvlM/Yf+B7IS3+lE8OhibxHfDUNwqEgsGQR5oapzpnQb/f8d0rZTGYRx0
XDPm2+SlW9KsWqTCr7A8vwBgo+uHOZLzmGp5/1tush8rPRSy3pFqy/8nckQIgqPNAB1kZRj6E1DY
19Jq5ofWiPmP1SXQ0VGFphFbpEdV51h47WKOHLMrG78N0e8cq4/hKDMtIlvzn9g2KCBfcJ5zvPOv
3X1dPhkhU/v/Hw1GPEulAmCBeX4eb4ZBkyZSchd+oWD4HAOz8PclQx3biabyczjm66K6C4T5qNo/
P0hz0cTmFMQpYvnnbsOTRscabqgEaLShTd73o1dr8QGwnIz59F67SMFrPqrnwsiAOf8tS5hOz7zu
JvBTSh2xJ3TL82a4GnWBN3pvoNnk2Wwz9vw8e5tgF3k2L45TU6Agu/OpRsI/HfZAYrjDBbCADlOV
jl9m3i6F6qIF2nz+4zrZj7Xo3uD6X5LDv/wQtK72STQkzVIZwuzBfm7ov/AncDlKvVjbHbpCIcn+
HM+8+esSl9nsEW/OpJ6fAU8V1OwLBQeZax3wsCXxQEG7qXh1kIbzOgt8AY+J2BYS/cWrbuGfoHdM
DnMrjAKcddgud79YC9LoEJFzfG/mYRj+5uBc5hHznhmrUJXXBGld3Rit1/lD9xI3dZMls+Kxz5BJ
t9JHmdL9cn0rsO8yFsBkeaPj9pkJU29ZJgFuO5CrbkmK8euEn7u7zcZfvjjL7ahPc+dDns+2B12t
DiTmgMe64mbR7/OC8+CXXjfuAfLtYgvUBNgNZtJyj7Dtaofsu3YLPndlRajp/kEVHa1qq20D4/1N
oCGmS8o1B4xG6jxiulhr1ho5BI4Hss5hM25Us0pNLoP8YO3Pm/Hup7FDZ7r3iYNuDMHeVHYBfxsC
NqOaXaqpzItYwJbMqUNBh2cNaLbrBbEicX6urT3yg5Zt4PLHullVCU7r3XO5+U9M7UbW6VxLizjb
mKW1eBs5ESwxiRvR9SfQSqhMHbZEvaKPKI43jedehlZW9EX8JLODv5SPtal9iPQr6/3ZxHMLEbZn
QxwMWH33cE0/ZLYQGPO8yk5wLpWw6cStIB5yVFz5O3fDN/wWeQAJaP4VdtEOUVav+j7m8+SVfjju
HiE8L0M2FKM1UFQ6/uEuJ92wsfxXe1wDD+DsmwwpCKVp1eQMpFRgFgn7KeJG36CgCrowDhz2ozD7
XfSmPlRY02fX4TdCgiZVvijaNhmozoWkqJua9voZntM+1ZS3nbLSbK76S2vDNoYXF8/+d29rpz8L
YxiXtbVgOj7Fb0vufd0NVuXvbirdyXSC41oqGX9n279e1lFNc2JAS2Xg1RrLSTK4qBFj8mmM0F4f
W0MubzLPB+4LiYosLg+7hYdyQt2gnUHvs9OCoZB2L37Ls9XqgxGeSeK2W5skgY+BU3h7PXEIuC95
iguk26jWNxBKixG7GhRaKSwSo0ihhbCUyYWlci/Ve/wM+pgK67cYWg1JmOzE6wR3DXRW6qrSNCfP
BLLyu8rDTUKMJjyjQi/Uv7RCUJ2DyCSEkDuc8Of9gqCmmW0jDOg48N7FFnbAgm9uMCmZRjUZO6sN
Ws1Zc0TJd/RJZrxsxM0c9dNm7Xnn0I1dJ3nAQiOJ0FMRi0qfGwbSIB4lotXw3Hx3jM1ZyziUlkyO
muQZtCDKhA3qOgMxt03oRfBXXMAB3Yr/NQnVgAPgykvbynFpAVNaqpfBWWX9tAC1fwYaUQKgfTw+
jF+5K75TDQPYsPiFTeQC8QP/ki8giqfjn4iKD0NPKxjPQkyJbAySUcB/TLAwnM8T8t9WYz5fi395
866xlcg6DDRMfkGazirC9yTFyduOVyOOCS7cgjZ1IJnOdDh35IySz5zvgqCm6nq+hlgdbIHeCmpI
XLg9NfTlvJyqwlv/i2LOASI1/EiNXp31QigpxbqRZ9m7uoyHzz83dsXRa7Z+L/n73r443pH1LBWq
t4mXc+PKyDcGrvY5e5k3OIAFHc5Op3XH7mFxO8xRLHLDVagTWH98uEagkTRQ3p3lyetSfvCAyVcD
zSh6Vt7tqAlkLjVADpX/iBgP2+3OUg5gxKzxRcmPLNUkLZXTjeDOgREwQYhrDsQv/TmZzEaWbMXz
mEGuRVXeKz5m285fBLNe0GDqadLQaIq8jMhiQL43TDQIVB94ncWDO+4pu+pmRMnwxQonv0cmz8cY
YIygY21oqYbLcx6BufCFHqlBvybiLjat2AmfbGVfNckzhZQiK42HXlkxvHCbjcbr92Athxmfn5nJ
ZzyG8cFlYW37PKnaSAY/qDpwC2M00yL/9HTab6TqCG+ED+feJQxZ+iKhm84OvHrAV1h0ybn3qhpp
ngpjVOPeiRbWJ3BZB2+F42cdE8DgAbq2LcKlQ13E/uAGtznmD3OqNRb9QJ6usLRJ/LbBpJbeWXKy
0X/hFcA4gisEtZRgNaDGMg9Xu99D87uGjKF0UhHR1qh9xqmOFYcqmTOcptF9aUz3SG94GNN8NcJs
sTL+TBOYMW2HIEaS0YWInTG9H6Uq82L0u/8V0dDoCF77IcstqDHE3MVn/WDq2bJvllZHKgM1+SXp
NAYU/ljulM/r/Um8u7LrAzU4ubclASsJBeC/v6AXDmKmU3eJNfJFMqyHUxy/xjcdq55Z4IQ2vJIS
e7IoMDvx0fOochmS2n7gzK7xvICoT/lOWc1rhC8ETLL26FcuI41PyVnGo1FnYSZYZPZWUuc8jvaT
TRCW7v1P/6dl8Fvrkh4XGs5oh5hLdlCj11/iien6B12+Oxrdt6YKaI3Y9aZ/XSRCKbmjQxDyo5wQ
6TPuBZmFTMyxFTPGv5/8G7hZDJS7oZxJMz4pqiHZvLXMFMJiFl5w7gNT+xnFV1C9prfCIagqSGZm
1F/6l7f/yHyXH3gwQWtMIHJhA/tqapF09dINv27c6yT0mK6K5o++Z0kX7brLRmxJ/yGWlbd0SB/z
WBKIX6tKaS6xj/LR5/4jHfNr8kWPRCUTUjmY8aGOfXjzXJBccdiYCpgMJtH3iFREQ6aTc4iWnkTV
xz5L8i3jynnC79d+7erRqElUf2Kb69sqIVMF/UW557IW3YSHB5hQ8D0RaWPcw712mkW7Mc/SFH9c
g+MpALdwCSqGh6DqYmlu923rlw4tsQCaloXAFpG4+W8OiH1VM1S4JFfd8T1+9EUDlDkeoy1YhTyT
cchssRrhnzCyD7PofrphBaYWHySFtlILvUzB9n+3WQ5gdgw6ZbUY0bCoFDu+GPCwI54YAbKjOOS0
79qA6+X9hIfqogpW0eKTfR5766EY5h+7BrlPki0Z2A62XDN1ilSKxtXiuZcqy5bewzbCNPCYvAUc
4AJHjVuVbv/sAUS4ZPMoWaXgAqXVao4Z5N/Ex0O1jYDicAW+oM/eZqcgBk+xf6jsi9v9JcO/38j+
Gu6kP6hXpVjnrv5aM6bgdJ/pYkeOyIFVzH4ORQleO+A3vDVNFNihmkF7PTjEe6J/iEdieQ7WO+u+
hYvBrn3QUo4mibBWl2FzynVPox3hR84BW8il4owfUV5HU5EyZ2kTyU+LkSSQu2sqxcLKDErsWIAr
ks7yPAL0JmABlMsojvuzimuSYr64vObMa6HiOiQqBS7Qo0qXWOGnm4uoJ6bs1rSrOYB/e24QHO9X
e14xwMW/L4VDMiOzRrtIjdzcfHdlWxAvwCvoMtlp1tdr0h2e4QM0hAXKYUnLBhehEVN5Uu4mWkbm
gtQA8tERw2VyQJBliGyjKFhWQ0NE1/h89BhC6WIeTVFbsYzzmCsax8bHvBK9UhRw7ldALLXYhydF
ivacih/dCeyza/C5A3nn9KuMYxNS9zmleL4+fKxMj3szv2hW0A/S/UnLnapHZt2EzAAyNSyAjOnM
+wXJO3Xq+sthnL25VH2DgjrPEsEmQNEAPeez7kdKLGTrUSA3TOwgxV6VXvX9r2Fv1jLyM1wFE2m4
5zdPXYoBXYDtz0Bd645pYj6E+KieCKLKfhkgvpAgLjDu9vDiJsDa1xhmgtAjBvT10j/uzDuHN9Ec
OchrjdNIGaYp5q2UzbOr15YBwFty69EWI0BZWcIalzZmWXcvuYsOpEtLIKl1HMLEMSUSxnoG9V7M
ndg4ZGY3QLKQcFzZwswMhmpuyg4CISTNXPsNeLCsGZRs943qDhYL0mCKC3okD56ZWhN3QLhCfi04
ChRyTufC3nN4cV/rImgPfZSeEfcXvp22y/dRRL+kHDXRi1m4o+O81llLQTMOM5dxu9JZNt0QPudI
jfNKrv6owS1iv2Ecb+WrNE7rwunevtoWWmiS9bPzQNOHf6w6WDaKwQioRE9/RNkfC4mwu/WUTq6v
kbGOAha909vaTemGM5Panu408vUdU7AfRaEkFEJ1WDeKet/aIhRdfa5c2rS3w9gwMuvJqaVOdEvu
M0ncHpaAYlOvTI0asgK3NyaL3AX7fv8TLBkSR5vlS7D+jxP9N2FRkcj7iKHrdaQGh7oqc54w+nMZ
0D/hTcqWM30TY3lUo1l/U5Udn18nZe4CZEe9SG+SmtaVPxXbS8ca231yOCuarZiVUK4HpPiqXvJT
VTid4btUztQ62athKRL3Tkg1tJFa1eo6Sh3rH6PJCAuYFXRWfjaTJeoJbb73yKmCKXPgesRp2g1l
fN20C86SE3xQVSAzUuVZNHjXH5xoYWhw45RVMc1bOMG3ajvr5y/LF+VYpIexb7NyBkBWpQ9j0Sqg
6FhP83Cd9wekrYdTBAGryyqx2uy4NXl2eCKczC0mXWbykqtSFJHy0ljJy/INZ/SNaUvh4LNVaE1Q
sZyRDoJjtLc/eDjYx0apX72YU+pm5s13wumD+wN/ZYXRx0m0st520oIjIgjEH+icK5bvuqtOrxKx
0lIXMcvKn6WWbG4UHCfw1cJ4GBEtYxR1fKM9hHhAXahlflvhu0omJ83Y6KKv/fEsLQiR+SgdsHAD
8LLz9RJnhRubazvYFiduyv5h50MwmTJ4VH8AGCWoELTuXH73RR4rGJ3yg9W7cG+W1nmpLXcKg15/
Tty8+Aty6UxTnXEd+NRcaec+H/wH0l9ffNRHJ/zXCx52uxSD8vQmQ25/6bCPImrfpI1LrHmALoEy
QMjX0lL+TBb3wkUdG1PybHzew7KHbYccZkHZOr1TPQhfdpDPQfnof4N4ZKXZDuua0patdNtpjf/l
KFG/fsr0/V4hYOHYO6Vo9P56CD4NhTOsJqAfyRsvkPimJ0boHGHknYIjUCzriF56EgTc9ALOQgs8
7FMQ4ib7La83gEc6gpT47JPt6ly1qa/GfRuHljVJYOr/7hKfLuwDtgfOI6OXL7v5rXhsOOIPDMwO
dKHqE8uquVTLVxOdc6SCzzTEKTS0I+7jDHOomnkSRPRQhdU+sXA9811h6L8fOlWXmhH1wam5GqDM
EXHg+BUF4wLZE+mvGw/D1inY3u2r1UcM82kCU9sAkSrbkiqcO8NoWOJPNU6Az7wWiU3lMtgwT8in
hDs532iZJuVnzhS+bWPUM5lmKnmFAgouYNzz8VlLnxopztEStgnDh1l33/iHO3e5x3DjbYppa+IR
+pgfxDIcSBNM1r2lUPm8S8wWgkhgsMxxG1L63s0tR2qLCa5kkHXIIGYfHjs3ZeFqN61YbzRIjgsU
Eif3vx/THF4F2DVCU5fY7ldX8yEthLeCnSUu64Ogf9HgCWwspw5UzXRaeiCWDWBGkBxL6NXbxgED
rUBIHjP+zakv4TOTZ85+lqAiK/pPIeLvim/nDDxvLGFv62K9yUZSkzPi2u1Dl3VSDj3yBwS85LDf
VEQTwdfUxuUQFYBxMG2N9s2oF5zgl4gEKxEVa5hb2hw8Gzrdy1ncA2+Tlc1iwjyVlH7LPC1jR3D2
e1LMJ/UaKdMMKNIZr/nZOczr1eiTvR42tUzse4qbnX1iljsY+yNAXvTQHA6kcIrRuCCkJgZAzbd2
xiCujYc+yQSNTbwT1ZeTrFrcluQNfY9r3VQXCrHRocgXe+RmpEKuRsOPqWhBsWtM4N3DkSojiN5s
WtRN7tstBRD7woo0v4eHkgN0FXXVDeTNcadhw/Wkl8lOUmtNSAkli+qF1lR0ZjJFcBVqPXiHEjin
9gRBC/VWefGx6r6jmGtHtGpDqeAJU5sY8/Y2BT2lI9AWA2sZ4NFB66cPmJz+37XBZ2MfQ20rQOFP
Q3HFsmGubTu6KOrCW/ud/JrQy2AGWll/58++SY6BheYn9dHjCKhnDrBEvcitRg+3v6Py+pry47Yr
jVRcShPGbJs1FLln5wBMLw4RKh2v+PP3DE+uyAWk3CmYqaq3+ZVGs6c2OAhgrAqA0VRPYVfqaKlr
mq/K9xcL3lkZVaIcIj2lEc/hsfqJ6mxBbIW+A4wOVlejBH5W/zpyYZmDCIaJRhBLvq+21oKKTZvC
1gGwAzRvlVMTIh2worwowfcuJg1OnyKHMSSl//XqValyu3/GI3fXIgQQtWzoWjSqCEgmftvvT5y3
g6ESEz7OZtYPxp+F5THexWiR+qDZLZjeJCcT8q7l5+FpuGD6T8dqrzBHOZlV/u1i7k6UJC2wqlr0
/1F+Glg7xn9c9BI1iHWduR4yu2EdDlI0WrtYzlcJ4ybiddLYtzKE7B4GC17fgne+kfO7ROZPG9KA
BeyOGKdAQ7P+1BBrdsgsvaPYGTwm6+ni8ZUouYyJILSx/HdVKt+83oAOYQOaBnQ3r05rKFEh8K1X
+/HYP8uSziZMVDRIZ0wBWfIao39OAU9RITQNG6oVJ4RotEg5DeqLjATE6yJkNMEYvPILIIvddOqf
AbGPxoptv5swwWdIeJ5+bd19VR+2FU8FkqwXS5Sg/+Xp3i5EU6E4YFOLwAJS1+3xPm4kaL3OoZMR
0bZrRVYdxBMqB/dn9KLc4aK+wl+w5syIcbaebL0PHy133G/VCgSqeZMmKSFbcbyPvFNazEKrSo52
ig9NuZKFlCqx88heO9bS5SLBy6C4hiu3lMLd06gQUZS4VQgV1pJBTJEDBdw5zGdO2ijxORE+1hK5
mvaV9OgsAdvCiaW44rXX3NKsv5AcqjT/KBr3ssy+p4uqa1kofC5PwXJaM9yx8MKPU17i3o2Ot0t3
5qGfJ1iPOmU2ct85u8LGrIc8AfVyQ11SeTnU7zk+96UmFJbRpETxFpUyVwtQCmts5kwpJ5475Y0k
YPnf5YCnE4fqz0uDb/bSkMbH0D9u9gawWxQkYC5V+gbwn0fa5+z76U9M3WIjrve+/QZf1r0nFBhy
vdyZyQInA3lXXx/APEpMlF/S5HpQ0dSqlDN9GVOZNiFEQmzSPMrmUPt52rnu9Mb57XD+bWvcbGj+
9sgK3GDMXhoANF/kq9d7pm/fUsu5xOzEHeQuzVIPzTtt3pfHK5nvVhUkzJKNYNQDQ/+CF7+HrldM
FtZQXHmydski+L9R/loj6Z9iwkAyzB4TMRuZ4OUcu9y/WBGvbL6O7hMRns1C2SvHBfRR6Ml8LeTy
NQsVQlqaJOzxOPWgZSMjOUong+ctZw+p5/VN6ahoDRZJVAFwbs6cKB+zow0E430aQy2rEZtV9Yq7
1pWngCMOeWVwRNNpQKgH4GxLceD6D17mZgRI8O0yCE8XsDFC2QVQh0S9pMqgKdfHHSsGzZYlSB/z
XDgzvPxpe068OVXFkPlBz/oSrjrvkdbVPfHb0GoSwdDQP8biTYFcmAMXokVVZwt9d6/9AeO63eiT
4BZljc6eKpFwzRAf935EnpBcEXVqCSOq3yBk+tBFSfDXjSW7FOPDSiTr+sXd6p2cbVgYUWQLka9o
U0ja2ml3mo3dS+FD/UU8S+dx6uqdLcW36gPWywvxBsAS2KZJyhC7YK7Gt48yk7PXIpA9tOS6TwKN
0e7aOLyUjeu7MverhTouwTXZIoY+LDHTFZJoOQFpoUCyd7BqiA4v07h1JmuYHqJ8Ra4KwF6IPwGM
i2UNkcn+buWWJaNJ5lP+fjuw7sgKf3c8Iea4rDCVpswOMrp4gpCBhaPfg04EgDQipc0LNopkYjzw
bgeasTI7PQlWZE8pnazaN9JCAciD1BxF9Fl3X5IvW4eWrOI8f7ipwsLt9QEvylMB44ZSoQQfp3di
zmeBZj2MWtblVpmoL9n+qFnMk2qEnpRtIqTW8zcqeu1zut9L1KkN/MyP6D0VmGx6bQmhx2aI7o+U
y9B0IhUBZageXkI1gLhaXRbby9W4KqaB/M+yOdaWXQczopcWPcHZVDTuDDzg+yJoaYM9rxKAIVGD
OXuTb6RbPFCPeobn0LJ3i95ZffCpoKTl1fO2AlD40XN5T+5QJzdf6YAouVN5k3McRBiR+HsTUad/
fmgHLypubKyWhufWnN0HZHyjFgqXZlSFqBCQbsBdGxC2/wyPKYr3Q14D0PNBoiDdsDB+ojxbu4fr
XX09VV85J6GAx8fGS6623Z0w84H79djmzpeC1E77auLxDlq+oCJDTeyH4hOXtIxa3DocfXZGky4B
nlh8sCmB7fw08xZey0uj/44TGU6KPqI1JvTzp/WTu+DFk7C9bgSEbFji4J26oXzDPFOKNUiWIDj5
AJtC1keNTcD7hsMxHj3cac/+IuC5b1R50xDruMbGai3b9iUKIq1vFdRERcuoSUt/B3EKix+4lqia
MVmsZd5Rhmi6xJs4XSZfjE3PzGT5iY0mDGbRZWZYol9D7VHc5bK8fVyruSuAmEX7Z4Ea1c0KneOg
nVEKll6inrKAOIN0zhYJbII9hf2wm2qjWtZtwYxqNJFogiIYgod2KZ6LvdUnA1Z1ePp5nfJQdfwV
H85EcyyDBSaTv1Bw5oXJMhf+eiLXap2xDVuIX0BOOmCamH5Iu3lflPRXYkop5MbG2c/8v55IqvAL
LPQflUCGvllyK3qp8F/Nemzl9Xej9LGfURyK/SC8DKuw5KdzzNmwhbNxPRsb4D2WgLlLAhS0TS+p
HOcPuq0h1W40P0YzHp6qZVcZmKGFht6qqym4r500Z9A08GdSwGOP+1M8w4iTGFfJPMXv+Xwghkey
iyAOSjDrVCRSD86YFSmmj2XLLEwbhz7pH3Q3ZWbi5YB30tgG0Cqi05Ws63G8mP4iZIwUyJG4S7Ho
9fK6p8cBR4I+5x8ZKYyRGqFPv/7GeGqLZCxGBQqlWr6OZOZA5jydbmJWcS9urNzIBEjUkh3YJGI0
vKL4iMZF4FNT5+CucZVHeU5xS76yk/vPnPyXIOj7gDJ0O+NIs81oQtrcqLF8mwe+ey+mMUAY9QUs
r5s2Itx2WP6b/BjCohoiEKxfSB7RCyOQz1OLUHhxOK2J+BSs6RpAYOevxO4D3CgB9MUlseMVQRwy
mCDSoBAwDNVPcLad/KdfSWI5o+CBox5se6nSfSBRr9+6jqn+VQRJoewkU0ht+RyRbyvyQ/5tLj0u
/Q0W0u0Dixid13Iu2u2s2u0v9aTJ2S+Ibv+DHGj4hpItwncqxUXOqBj80YSi6KbPuC4sqMastFNy
iXAYyWCS3lboieaRJly8s83V+27J+sWR5c5i8YjunAKblMtrEo0jIJ3nvQBOwxLcn72A0tSL3g+w
YVgPNZtzdV7JWjG0ihRGbHpZmVQ+UFvGmUizQ9kjV/vEqInwrmAXR2gqZZ3v7MzSHmzNdWZht7l8
rHV6WsxxHliqOwi5+aBJEffnk2a6IP6mPk/azdCyCK9YPx9F31PgjeKVt63OLuLX/tERFSc7gxA4
BU16PpMnf+9k14H9Ot00xtWwzAapL5d7Z2xQOaGKnJuQX/z8vTsBFbPaQ0YO0L0v9Ph+T0oEsxtC
bNtvW5AV36M2KtRmfJ1YkQgIP4Y9BTN0Q5qlmNfybKspqc4nI2X4bBToRGjS781fztD5cru1Yw4X
u7q8b9GLPvkGNbcpqRKMrfODcAteDsGS3V30W+C9fOe+VKZ662KCu2lUn2V4nJ6oFFNr1EyHFLdq
niJ3HF1aiVG5xWGg0ibw8u/aX7jIF+Lel6Fd71elX3Svq8UqxXlzcdo40vYHt0WSSLyvK/rgra/t
A+/rV3d7HgoC7GNCxE2IIySr2ejmwW7pH9T1q/vASOxrnJQ1jnubH2buWhvdkiPWUjMFa4dWO9CK
rhzuvrtUGyGmZJbjny320/8YePM95N6IXDbUvnLag7PgcarWJYO1rXIHnif0EBXTAD3GZwKs5lk3
suf/p0B22S8QI+UXEzpBoPXUrWRL+xJxVUhbfVU6XEs2jGRYBZkoj6GLeVx9BJHrW3KbBISscnXb
7DiTswGdmc4xVjb3RyUSmk4+rYf3TLZ9daNW3B7wR/SZ5nxqrvL6yGhKtN2GgdF/Pt/0kP6+l46a
Eilfbpk6e7llTxke8GSIV6bDHYODK6Jn5mEL2AmwLEenIraWjZkxm2YxomVH+BmHZLZIWFLuo2UL
prOqiF7QirB2VoyrHhcCg+qmSg6YLfnwGLKxbYdv2t86Bkl/sLxEDePr4y1/4U9Y8RD9BxteCl+N
vc63bhWGs95pbutI1ZeTaxJQxw7HlBHdB/LP4WbrdypHwh73HAeaLshMgFNcIgDg1ndSvHcRKWf4
NeiaZdgOaHU9i77dG0pJ4UrhPF4ykTkbPyzcfC4WtcyELslq7GofO11RKiGhe3Ilx8WTaCeP72hR
61+mGRtbs8bNVrlAOw9PGQtwshGD5BHezT1nXB/A2jpYImzus7WhbDyumhKV+vOamqoB0BjosjT5
CH3IITXf3FVvonXXNtQ7Yo07r/yjMgwXts46YDDwsGvw2CkLCKMWw3s6q79jG+bzyZC3Uxg5mR1s
94xTWCxvkuoruGR10dH8hzGQYvuEXhWzhBIyuCSOdLtASB1XciMlkH5Gd8y4BlhLFHi7PWHgA8zt
bgLHq4ierE3WEoXQ25x4GbcmswOwbZd38p+i8kmVVO9saEZcN7cSNSZyxdkIFaVwVAvyayM7cE4X
PY/IRmXY1XBTlHuzQBN/8wS3NDPHtFdFBM262TztI2FxHnsbl5gHj58qYZ/kHNRkzJLO4Qb4JBk2
fMDSLttiSRs/w6Xpx3Sdv0WOZVcZlAIkq1OI4Qy4p3ElustOuMXkFmOUktnVxy4+54yL/eZltaeK
7kSLDaiSKTGFs0zrZDl6p9nP6MkeSyv1cJOogdIlhPfTK/gkRXvb5JTDwFY5H9JbHtw387ZvHibd
k70jWfru7NNIqVmZjQn1WN5+2DsYn7gnyu9v5Y+U81ZTA2JXCpvquIGyAQPp2TwOaHgk2D6BcGg2
vvc4cPGS7UP6PgzK0q1RnBy2oQ4x5zUOvSa2CDJqASSJzlDm/v/Md+yy6URaofKQbzC1aTlUD5e5
hV2CCDY0bKh6XTRz0PauXMaQCO+nWatvt31kNfOAgVNq0TM2Hvu4WdkwBXd+F3HFEvEB7hexezvO
rTd+5CLh4Uu98FkU8xsFNHohdIytebM35IcXIkfy+F/hA/qOFTv9jZgE+9khIrkFN674P1YS261x
O2RJBwOVdYIgz+aU80te4LuaFGte0SMwoqC/EtkPYS6y4VelbQcuFiwT4DZa7yuzAqtZSWPd0e10
vDxnfAgWZandNTAKnXPCJC0PlL1net7llGQNzS4rVreN/sBNq0ZpBG8Ocx3+zTxLAjkGb2dGBKsR
aKwkGdc0r91PBEpGBDKdQZX1u/ObxTgDi0KEtV4vzF695z25QDNgXDX1l4E/r7re1QrVzf4t5ky2
8sq1btisLPvVceHClYiedNVU6gFTX8srLDXBzgXSiyTlLdtIwRQguR7754QIXTs96v7I5aR2WMQ8
Bao5m7H0jM/NGCm2aXo8ZMuL9IgZVUChlmvjWznqU1vB1mhM/HDd3Xvavtg0/vWBj7CpZGHYwkYW
1pEeC6e8dYDMq0kzyz6uqgASQzd7HCjA9BlSAeNLoGaqkbI0zGHTG1OpVNmiZfEQsPFcR75rvXqN
Q4vEl3LD5rzyxmufU7P/NsM1Aszux1C/egaLQFBew0XBtxzJlMpW0sxoiJ3eYTcer6wupfm2poo1
vO+9a6vM+YbDR+8vckuJimCcRLIBHWQlzXINAsnwzxb50DQmtz32lxzLaSym0YnuFR7w/wZnk32C
Poa6CEjBkzYCQxjl0Ga1gyOKnR42BuULg+OnOjPLytdYl0cV4d5EmpyrS/Hm4f5BK5fkaxaU6Efu
WU1g8GnBEJ3fVJon5EIri7cnMLH8+heBVSo6maGVUPgrn4s3hKtNzbV75HoihfVc1M9YNTA7c3Sm
0HgvkCFxdyPedx3QnQcCqPw0YqjghND2nVvqXQATl6T+RwkEf9I4j1917P+OCB3iUE/HJnvt0Cph
XReFDXyFgt6ASbaS5vsRDE0G0XcKP6e4taiY4js1z8WE7SHtuNEckU2+E3axfsx1D1nqXHNDT5XB
PV+VVf+iYKsQNFBe/c5AL9cdUrBfOMU1UO6kE2EZtGKAiQ6VCk19SuAuFdPA6WtUSF7xZ7Ut/dPz
nUkBpkGWQRMJJNmXThQkCDxR9BCDrldcTZxPoGC1cyIiyb0gRq79V396dPpZTp78ffF6XXBHvrIy
x2hB4nqod5uC2tsi8kOAOzGYZAm8keuJcbUcYL8zzL+4cs6M4+Hgd0JUQse+9T6C048TAhnRyiKr
xowyXfAJ9nm69qww1o9knl2oeWTljzNGsLoHiHtofWLOD3FscyYXvfojqc98OeSxBh/Mtxhptelx
kfdMiGXUPi1Z6oOunPJrZh/i71neQGN4hoswLJmzdVjnDxhYswQ2i2pc6ubojGh6t34ktKKgQZzO
2vDTtbV+5DuDTXXCUW+YKTur+2BPfHv/v1DMkLMaNdeHXyk0ipMh/IYuaYRpLm7QHo2tXDk1LhI9
uEFQL/5JTr0ZED3CSkGdihV3DSKrCQ7iFSA5NMV/NxF/oA5gpUajGTfGl2DrrrnxaIbX9RpB0Qz3
pOp7gnsC7mJNMeybEIjnefiEtqCNyTBm0KqlK8xuaU6ujs6eEypcjFQaxZp/ADtT/Ytw5gmM+YRH
EoZTxjLrbT19GTUSLFrZz9aSMqQg9tc3tr8Tow4iZ4rwJ5ou/ToewZd3PMYfcJp6O60CMRwzGOpM
C6zXXv2+yGOmhw9rjtS+j42/Ep0CKqgYJLn2w/WLibtlr2+uiJijZvivlL7oM2fuY4bCqhPhZWDE
/WzrKehXzuK7DcjhH++YPm4BFLpvK1C3VOcvX4Cbo+YwgL5mnWtanpSNFVGqMlgNM7I4x+d5xUn8
FcxB45COPbE7MbZpnkISIQPBYSbVbwzOKoXXpBz8JjgTY8IsKnnqIz1j08cPWe8FlocX2zDidE2c
5R7F4P4Xukcw4JNUnhgzq8FGLcBLF0VrMpODGYARZpjHh6WlDSf5bjHKrrDW42pQODEbFVl94kna
s/WtzO7kBgvpsQO5/8o9COIYTc2tqoYfevA4q3SwaXxjAQ4nDJPQHNaNAbPSSmie3y669hklwbtH
6p+NEsQ1pYqRDlg1USgecig1RSwsbcvOGQ5TgcdOeIm7kWI6VBRWxeXatXfzNVCEvCstPvAUaF6l
aYASndZZfJEWsSDdf9I8Bzw5I7Jx1rtzPEUxPVG51ZZz7bEtBR+7sEMLFuVJQNNljzi7tg6dCu8E
KUvnUIBCYiFLsiuVVw2IE7ExHvTF92+GQ1V2Oc/7B18CXTZQcYpD+la6IrKN8O/l2txOHeIvFHCZ
2XpBojU5jbzKCTTnWp9Kl9S1Hb0xcYkVrifYph+P5mScnJYvGF1qrbZR/NwTgIbRlIZuLDvYj2so
MmBce9tkUXRnc7Gu861l9q/TvOuskaNso2qA3zT5R9qmK3/UCCaLfQ++oa3qwhqyVvsdKE1g0Vw9
r3Xy926MZOoFf16l2AzqOnf3N0WjUfgiaMaTl0t8gBUfG893fsOsz1HaYwWfCIZEVmOLJl5z76cT
g7IZNBhYpulY2Ke0Brgq2xnNSzet0sZAvQMvwtyrsE2DapG1m8mqlwPEDi8rcxj1cUZk6nysqMB3
SMK5v54OvwcI3K+/ADLHB9DAwB55Myh2USfiy1E1d92LlX2Hq4VGrnGfwslUCoSk1Xl7/AUaVZvW
bEx2JAEW8OJpR1UaLskyOyhDWNCg298kAE9bPjba6a0FF418XdLtJjwVcU2Jb5y0EOmDtyAzDr/r
L7Z2MENqWCbPIAXQmIlYH3BFjKhFz/kt7qqrv1JP7JGFdu7bt3XN2irf7JLASIxO7DgAlDELYbaP
zU+oTAthneT0MBZDek5fC8HDtLlv9oiMwwnwlrdVCI92C547A+Wo/sgokx2aelDNoP9AbVzGlYiy
INTNAPBgDBT5cY+jhuDrk5PUlTSNbTMLmI4jODoOib4GUNsKpAvY2Jh3ePI9DLRuaTyMkYcW7ufp
jGaxoabt7UfzS+x8cGjaBuzHfcxq16gxeXYXAvC9PKaGz1hSj1juomDXce2/1Pq2c91U5JlVULlO
eenc3EArDwBQXpZEfeni9ClroaUd2AtVYbP9cacJQlko3u8o4YNPIcE0uelptv0k+0Zsx5CUFH5+
yghrsBu0iQeus1r8MTGw/iSgAJGd4XZ2oCoPzp+tm37VWdLfgvzBPss6Wsn8/Dfj+n/YSCG7aoyT
BZsPaUrrKzMmBDFJUjETrOMXaJudUTUvwMDiC+rPglyX/dvbQeNH55j2uwoXgzpNv318EqRuEKof
HuxQ6WWkyzefqukT1J4IKmMJyJemjZf6RLhHUbq1RV1WBkSlUxH6Ke6lQAwv2pFQmUd/86nQlfPh
jvtbQATomX1PbGKNuXYotJvu31Qc9kj9Z6/XW2q1Lsy3EiW7yn6c28AAZLfdtyrr2x+cumJWi9eK
DP5GhgdCBLDnuHmQowPinRLwAY2Y5EYDpFirfF3QUl4D6d9TfYa6YPtwG76Ghwuaw7Upq8Mys7uU
LjfIwOPvD/sw03u8LOYyEhytGyF8Gr6iw4G41OeG9/+lFZQVBTUEm1T7ilC2bDlXfcdFKncTp5cW
zUtS3v75n/gpkdl2LEU6oluUhHIk/pEvSSPgmxu1R0SNh8WusOg0f15U5yKvb/DkgO6npU/2DAuC
oaKIuuvJfguW7FxhyQ+h5pxg1/2+lG6AT0yf54/KImwGMfsQwldcOcVTDVyP/vQjiEx/SqABKEXz
rbWUk8QgybjFfKruhxaRI18DLm8eYa2QDs0rNTJWZXZkzO/UeVBKeX90Ppx3Nk/J36ATZEQM0Ivl
6I9yHx+tPDDbtLpLh+2YOVCItdhonuDEUtmBPtV0vG22/WKf2bQohTzmyCax7vRlYW6S8iBgoXaL
YLG5qPn+v5vYALqFf+HRxuDucvaUSQ0lHKzHcFLH+WMXh//GC+TCoMWK2HjBCqAThYiONbKrwG6c
14qg5tNUdoMfq3fMf/XJ7rWoUZbsHWV1A3mOQzTkZxkJLDnq8/E3yFtM8GD3hdQ+8Jflgs4GSE4v
0mbosxcWd7st409zj7rTDj9kPnz68DbGvM/FSrefzShsq3Yypt8N0RR1r6R4DKzOp0Bk1fmDwqUr
h3y6Ac5/icTfI/OiGqK9PuEno2drEGxZ7b/6cjqijsEypM22VN8wSl0A+41cr8Z7/3imfbSTiNtb
VVrJJ7KrHrvpsszmi9f4lNqKBpopB87B5Rwb6MTo27G4tT4RLzU5hdARjBYhiIn5MRFO4+u4aFgW
DHAehBoW/w17Irrs+U7AbQNMqzB0/2HGap0rGg59S/VUz7yv+5+IZjd384V6H2RoVQVkVQm3yGx6
lr8QEVXNzmsVNkzUSmmwbAoP2kBloxvMbfLbG3DscD/tuGoz5Pl6owT0GJus2h73gI3+MLHVdZl4
8xKgEzeyc8N9d7W46yTFqoljhFk+VzS3rr9PXvZgOdqsmkiazv0A3+/GmJEovsNk7zYRduRPU6dy
/GZ9zXUNP6gFw8nDRcefJEHLTnA+F5dQCpNC5xKw0ttlfsuMIIQ+IXYbHMZNRlOv+oepkuhWbWFx
jcBCzSbbivYv3folJPxC8v4Api5KtHwjn4z9qNxue8/3b+T6f56YmfH5OFZjANwQE8+MWfxmZmAu
k60NXpRd1JtR3OEP6A2a4XbnYcqrLs7rlsGEmbT3wDc+4hOVpOb0jzmieklC0bySA97FuZhF3bPR
og7+QOug5ct6Vez+ELS8AHnnSuvY5fHX16t983lg+ZdInx9APyYJBbMmA1M2bLWT1Cj1cShCtK/u
A88lFOp+nUGtJVMuh9k2RV+4ShXNmPB2499jUr9VtJhy5W4cMh5POCHvq1VSAsXMQy2Jx98pT3V0
syH7NhpO13QIwyYujmKOVeSKWJoBsZ+UAV8cFEI3I7DjEGmDQ0wDInKGjpftwFCjcblqt8Aa/8RI
kYsqqVcvA2++A/R8uHVZEcMm7R8dPuxyWfTV+7ZkJiSoHZvdCs89m0rzW0vpNfrdXbyC9APUPiRZ
uM4R1OZnYF8J8BSqcM5g5AUAP+xQ09CYELHL6emOrwYxIbHDcHw2Feu1IENuh7xlvhBSs7QqdTGW
OaeD1s56DIRrhcdX0fqPsIv5kgm+IA+3L8Al22waQ79WDgUT3/IvfnBe4KspJvbvl5SRqS3krmbt
FjH9jZv7BK2zqUoF9Cbwi86NmHa3IgyVvy/QA3aTCWrVQJQqRt3ByiQlCi0uSkZFNapx8uychcG7
LTNtdCV22sxXdfzvI0/xB272CMlleI4Fq9xwsYn6shIUBKrKgQMHUGX4++fX1ADxDIihB+DC3qe/
iWq5zbrq0NmUN7qaRxcvHdnee5wxRU9KCBDzEyUaYLlpXkRQut4+tVBU9FXbx2KKXVBj7eCxwutt
WdO4yXcCnbwjuWesz8/iikyzJNwRONQPCXawHZL1Iq3jiuDO+x4NpZ/T57dcTP71BehNNrW7T4Oi
/BbfcTx2Yl7O5YHejPG52gzH7FGTibjSWvrza9/I9Bo20/WTgE12Swf1LpiNtfntkR6UgppS4aYT
jnTd+Mjs2VkWppe54y25Z8ZMcwQrECQ+PaNoAp4AGFiz30IzA6Sts2j2NQCbtJa7icnc4ddEMa5a
FkKOptQ27kPcX2KJXInv9skGL1KUDhKKIi+qOfk30UFVqFm3wGumvgHio8ZRhp96eGP2CGvSAwsL
qM0pQaydvp1csyilsEG2yoohmqGP8WpsTecCUIuYgXWN10qB3NzBtfyw6Ift8CJxLm/OjRFVJ2Yh
MUSq/VZYuxrKtWyUtfT2RBkkzXhTb/i74EnSv0o25/X7JLec9nGPAkv8svUYDgSnvixeUklW1v1U
S+JJy4P4J76fTxkMJGuCTqD1Gu1eHlYQQYhhwYu5SDNqzxX9VBJL3bMAWpwKeNaXsgK/Pnqf3+YS
v24OX0OxzES00qmpl7RARZ9u2HqeEaMnF+gg35Ag4CeZp2oZG1j8oxV4UUStcqrz4tX5kJ+U5+Mk
6e4SqW5EbuOG2I8WA/5agebgiwrpJJiobFY5l4cGVtOot5SsKG2/HgR5Xf8E83lBoghsJGNZXY6S
kp55LLK/waUthcuXz3xtUm2w9c7auWIozn+jFJOuVGnLOoIQBF3U0jfB0s36BNzAWSAwrR+t9S9X
EAxqHjhX7KAKBc64AEYlI/A5BAM5d5Luvh11Qnm2tgAkeV5nKCnUShQXz/35FBZ2uvSqAZUe51p1
Rm2UzStgh0Po37ht352Rfw0tz/LZD7htoxbKbpjbuzTKwmkR5W89uQu6wAx90YMLf/XV6rBBSJ2S
O1Ycn1TcJM3rWm46r4GI38JLc43pfallx+P0liUpIgftGmZXHIeX64LQfD7jtM3DO7poCaWECYju
u3Obuz5qn6ikJuK8u0thjf9zxpuX8dFHucESaJr6NlJQjGqk1lL49sKYdQ5BZ+dIaUt+Uqv8cecQ
hEaYyA8PHPQBkGJzRdr1MYLaJ9xlFEu+I4yoIPdLzzZJ0TFBZ6pwfRzT52HQCBcfSQeKEto9NKFA
Vb9t4Nvzdl5O2u3Q9uf2GE6ha04khV9k2+0kKd+vR8tYpMaZt5P0XSKqsEE3jDGEJ3Ryz/pBSJVk
lQHBWVCMl06LpZv6FHHnrqJhX5lID4EGRjMlt3CkuIvJt/VCI82nDnMhIZuOXDN4rR1KdYnnpOuu
HHakg+HijKUtAGruLUpxlIR9PfDqot+wTFSVumoQy+/uQGBH+e3N+KMVqnFhlcxcYRT8ulu0Pdj0
9IPuxpgV7hx4fDvNKsTeLfM9d21Ylr/3lhIL5EzyHRzIcyN8u0TLCwBeekWHW0t0nKCPAvSJBYmv
VPy9TBnbV//3XScl60CqjZbfeSrVsZILxRLdQpzeQOcf7yUxO5TMcgildFe48fT7ECHMmP//qhTk
ikdFb2dbuS7qrImnKoXi9xznq+7g7EJFwTNZ5XtTUJJ+esaSsgzV0YhGJHlGlQWA7ytuPCYsJu0S
IpvE65Mra7GeNMhct7FrgH5wMi4OWMcllNA+yL77Bk5PG0qavoTcDK4PPFzck7W/yxsMW6J6cfdW
aJR7v+8g3Y5JiJS5+lYwat9LGr0jUl4nO3LaVTCXCjVtIM5r0FjCm69Rz14Kt/mNzZ3wN0a0CMHl
yTNsLf1oWIN/rjhO4sUP+zc8BGZEHWv65ig1bN1jKCcGlexFgjgUW4GlJ5qyZJZ00EFo4ohMwMq2
FAII1oWsdIUFFgSV/YD0TXOiIZrCW2g+IK4fVyDvMwOq8kMfS+drI6S8fyZBun72MR5Ra9BcN6NF
CrK3UuB9pqk1MjbXZtUb68d4/xFbZpNa3pBnIzX2xwPp4VLSrLnZn2T6d7bcPqYRIStSieOKZpqg
5kWYnwdokkfHFqi1uKiKDVwvWRqIWVJPgR9p/jWQ/xgouLNfP9bFTOzNpaM+pSkWdlLvD1ixr0F3
jBQU1ES0AkCI4B4x0NTdlo1rIXQSyV8wLf8fBlrg7tLmHe55YO57haaphVp3dU3esgDquD5+lgsp
sMBnPD7X+FUkSyGomltUcWLImyJM3wyMd51Eka5UnOHCENilAQUNNJC1K0AWEvRybv0JaYamx4p4
6/dyyfHR/4Z83FbP08tnQji42bPjdBrAql7SwWZqycm5qBAs8r5bE+H0yA+SL9OVhrpEIiTRdvbe
dIZa9yeNrRbZxb8nVYPE7KuFjbu+/stsrTIN+HFNhG94S1DtK9jIAlFM8p+l2pfylfpSRHeON1Dh
drqCxdLn5mbCkvySu3TLplNfQJcyIgKNc9DfU6z7yjwpr8gywOnC5B2hBSBZRjgh+rKeow2ZoNUS
5qEYn5zen2G+aICE3LZIuH8lzBitTTuQfuRofZ3sXFtUhvzaPyQBBVtEFBdKH0Ykq+yzgH9w18Jj
SZzXG4s4zmDEuBVwO1ltKw/oX66tWuM9rp9Wgu/8Is4iEl1KFVszLTNRdeCoWr//rxFufynyKeda
BJPgzZ3f765J8jkCXu7mPPaPupkce4RfPYcugaF1iikKRJwJbSpxMtQkuwnzBtNsAQuCzX3+xt1M
X2vR0bjf4GW80YvOekoJpR9yfFgAbnmuCuPWsaiB/YltK/81Y+zzGO/rtHJ+64AqHI031cricmY/
ak0yxCLIUOYvb8oeC/TrUNIvLcqD1FJMaxP6LALqHKPZckLJi01ZrgrGiZQruGy/DpyuI/MAiWy0
bMFFtZNJtB1CloYxdBUn8p7tB1bM8utFxMWbIWE1rTX0n7sP4B2wfMeSIx3oVFNzhDy3PNqo9pQ4
cxHnBJo74y2ZKy0QNXFwSxc5RNPNoMQZbE7xS4wlXj9cfEVjdl1B4KQRzUdJ2OkxwDmEDFk9mI9x
v3UtYnnUNv/66wG6jEaLGHb49z/sN6NTDXIq+Qop/eOamo/v/F84Ywuudmxsl1GqCYSE/oY4zJ6E
mMf7FvEoJj6IDFOb+o7UpIfg4SP0LoYxI0V/Ee2cmThbtKKWacRiUAS8W8I/5DCLPr6yEDIJhvyo
nGqfnPBLOaYMgZLAo9VsD1ogOnnQIqT8gHjtmTTfYwAHaz55ib9+T3X49GnsKzfOvonSCqzHe+Z6
tUFFdCjDjWwPUq6Nh3DhrtgoLp0USKhK0NElumRNqLDpkzVagE/2wV+mcCzG2VgzAk6eOalMiD9n
YKoJv9mPXZtvpk3vajzd4fU6GpXmNjSX1ob1YoavFpuvjXsRlHgOrM5+zMOBAkCupEDkrlU1J6Od
uOMYrU6a5m4mcL266PQjhq2L+p5ZfOAhL4mEKaCBNv507MzvFUUYLHx5wQ+FSGya5hylzFFmEusx
hVnAUhWofRagItJKMlJCMZqPToRZruu9ZYcxmjZYAviB5sca+mQdU9Aj6hbQw/voVAlMRV7OBVe6
9YdeD3RnK7pE8w6ICElKQmDKNVZ5SvBLDN5wcTIV+XGNH9IU7uiK2fclxv5wr1UM04UIKHpMAfyM
t7UqPtUbRu17oGFun1rI4aH9IGByG0hzwU8lHTmnOF1lYHLT2/dZKwK+ucA7Y3F5xHW1TRBMfTq4
1cJWoci6O4bmmhxPDHFtkWnbvYUB90mwjdA9SIxjOlwsiBH+32dgOzd0wHmbnkwAWcT9R7vmPdt4
421UUl5bAvQTzPvLKW9pfB353h3HOmAG1IFDZvbXioah/rGkmeNNzsAcAk/AMtJmLz/kH1e+IdrD
ApBTiMxDjwPgt2Ie0HrYX3fIPQzdj/hioqWyvAHMyVwITDwhhJOYtBj970qpHIrE90oAanqEFZNC
BCOTwfzrWJVFjkPvigWK2eQvyOppoGjMo+R2kjoMKG6Koh3TFZwWFznSUwGCJzsZpXy9SQQ1azJ2
+qvUL5YErUyRC/JIPFOC/wdJBSTj+ajEfTuWFM3D8/IRo29ZbtvOzs1I3Po/iyJ2yDmITBx9nIcb
oSmJ4/9j5+iovpMUB1qvU22qHCX7jGWAe5FKBg/wK7KeaSGqjAq2L6bqsTfCkEWEWWaWvLZz+ztv
+VwStb1bsVOr4L0N+sIMmAmLnZYcI03faHIMMlC/TuG7F81HXrGBiPQJ4RoUqJaZzlE3CfYh1szW
YeN94HC0v6uV7PWC1owduPypSkkzd3wSaJChCYcEldZem1YgnHEPnJ5ZMRSVmfy9ZDw1KI9q08HM
DSNru2ye0YF5Dm8Tqr14F3QGAGDk93RPYB49k+hTF2iQdqkLSEAC9kIPOcooIYpitRMXUrckI6Y1
2Y5ILcKkSrUWWsd7GFE7cbqTyFdUI8SO3RV0Oy571Ik0nM/1BXMPFr/38pWWqkHVOjdQvzVMidJF
lQQJ0sJLp7BDcQbC1PheYWi9V54zU8SRgS9Ss7KPP3b/50v90fk1ydT/GegD6YHeFsMc1YzsKp3B
PLvI4gAm0Sw1hVfZoknPn+kqS8tg3p3nKkeS4mh002RY18Q89SbfE0eMO+/FeCdfI+kYWr+RMeBt
PsU6VDkdp7tr3cE9SjOFDHOLIt8fHkJjccR8uXmd59DevMZkKgLAdhyqoXDi9psJvHQTzZuId87P
AsCCNFW6vWbPGXa9ljk6JYM3xrr3C0jiUS68JqYkefmFugkue39IYgZYUVaq27T+PHyP9lE8K2NA
YcEOFK/+6SJH2D3/qEVf40MNVpW8rMEzkGFwqvGOQ+HK7DG75eBxjKQGnKK39+BXS8erI/L9MzsF
wlD57OLhlngfIsXwLWgXRVbcztLrJzg4ZkM5wb1qkxQE05n2txyZ59XQoDFd4eiXikl1uAMWLWzt
gBmulrb5CR7akWIMdDzU/29cm/inGK9N69Td1WFnlBr+fU8tsED3+lEBG/sVomtSmne+QxtyFGeM
ofhfoC0rk5Ms1H9L42BpNS1f/tTbpx4xHUlKyw9jQxm5vCKrdm0ZIC7ZchfywjvB4+vyLpH45WUD
m047zR4lmtgm52TfOlgNSbr+nJvbPLgJhyKvT6rgUO5gFONQ1r0T99iahszdS4hzDcsjKmfKL08w
PT5IevkI2n5bc3bIO1IKNxLx2bLJz4Za6sjG6+rjgdmj/RFyUIPbnvCFIV/WU4fLOY0jZNvNG9bS
htUr0nzL+0YXCCKj8XFfzPmWndN9ebaZ6DOje7mmPyCp/yL9UHQJl4O97YoZf/DPYX2Q6YhUluxN
8oQG8iyaTckOLMIKSBNce/xn77R9i+ZEMlnFyl66abvpgy0LmYSENHhjz15p5gURcwVnYhmWeGPD
Y1dO/NgFemkCz+rjCzsWdu+1nNdXSnW5kFogpgnK/yPtlqMPBFAWwQ/yMFtqgAURmyzqUQpOBCPM
YvHVS8q3766iAgEUpMA9gnzY5GucbKE6waoeCKnmJPsSazVtHK7P6s/9EdEtn5AgHfbAowkZcK87
QrdR80IDe3Gba/PBZtQ03KvmPFAGcA79100CdbyKevmfrFPI0L2UDKsG2QdqNxzOLRHkHVHUbR8C
t2ga9VSlJjK7IB09LDr94jI1fSs9+8XMOJPH8zMcboFyvh7ugOzdk1wILRJiIc9Gic8o2HYefSiB
CFjsAYEY6Oq0ubneN+Hj34ap+YG/XiQLr5rGhvTsJiZ9PvUgDepn/Q5xwDnM40YwtdkGYlRLUL//
/3HwDA5ufx4TnMhslRoyXm4VDh+Onng/uiAsrPsxjVD6JplYkDMG6ZT6cQn59HBMMrrc6ed2HG1t
uQdg8Zenir5wXFiHMOQKEdp5AbkRvx/OiYw0Jf7rGXV3lM7ZFOrSk7P/Q0yoFrjjtngP8Ujadbs8
SD0nt7ZruoJ+7Pg9vSKjfBWDnaXm5aLBHIzQkOTPZDBQic4pN4h3/uofytd54cEe+2FEFXq96D+l
cDFtxKRRE46WWDc8yoY08qAISoIXmJLRi+lNzU1yTWR68D49rCYQLlORm5TqmiGjA+rDyUcB+00E
0pXCqPdjS8Lft7vQr7wb3mgFoOu1k+wsVDJb8tWofDrTS+XO8nWjKDP0N0vFnF97Nz2OhKOzDPlf
9acDDuCSikaRVsKIVocg8BPXmVZy2dzMYCqspH112EQrKL4PJZIX21rwuNtR4EgwNI8he5uRwn0R
ItpzM6Jj5JaCoTWNq3pUrNTvhGlT0WDWMqO2EElRirVjye03OasQHzs01SjDGCRJls0yimGXBelQ
I7PIKcm/jS3TlVUYCPJ2hKSu23qmTPFAhUU5n9sM7wRvUwo4921LA4hKJ0mqEU4H81UD0IdjPduk
3wnBtK1CyobazCo0MF7CTIyW8prWSw5CH342ekH1W3R94lM7GafBuswvtrzJFsOA+MGymTyf1BcI
MUPSNGwn+6Dn0xpc8/wrFkjn9qkuvuHZEckZChrnaA6rZ3dGvMIcFYgsjEeAHe2rSbQ5h7Hxz2yu
6W1JPgLAymRwhxOI+YygpErgUzlr/t6q4aFOMrWYzAWi5o3wPHkNXeSBsarcD2qn2U/NeFydZCXy
t7eftI4PAWX4nMv4/X2TvE9g1ZrbWdtK4wiBeQFV0wh12+OejAeFIQlVgXhzY1BQjpRBMIkobNqs
fhKXadT14Rnvr+xTOcXItCC5T49flp6k1OxPLghFgTGnIoCU04vY69eBCFMv7HVjO9muBnDu7Hlq
+2P/90LJsbyDvydQ4rV7qXPLGysvj/UMyZr82RVTtDaf9KTX8ij4v7UJxkLlIgsF6HjBIDyptImA
a32eNIwH6FrvDw2Kz1/GlHDKSl5zN1P5bpKB2/UQP5YXbB5mLhik6YIlsb8i01DnImfJtc358mDN
B8EheJTooKSBcrTKJNE2iDFl9jg2trfocl8MXe5tXaTf+3gBggPLjqtIZxyM4OFcd5K9c+N1584y
xSSLOdD/Zr/v7vILVPF5C4nWIYNkn6cHOCTjKz9f/dinv3oOSdq9u6qUzXzRnVlH9faaE1mdmvvL
yWbcPV01rQJtpPn/OLgxv4mQdcjIVo1G6u5KT+IXeoztqr1cvAlw7kfKmeM/aE4g20uCj6Cb0Yrz
sm1S6R3kOpzd4Q/dtL4ZT0/eXQnrGFOKDt1XXudbwoAvnqsmf7iwnVYTV7YfDX030vlNc8/k9dZM
iQ4l+OCaZteS9w8MBlqn12jRAYowj5UIBcxAp+Oz1gUJphoP3gIGuCITp6ytOrdP5ikrUd2pW52h
ghMfyi4NhN0uvFIhyQw69UBAf5dvJm35v7rdIYdaipdihbkX1UpbdYldtSbAMx4j8icIQxg+5vyx
3DybtB2svIqkYNlIKf04hcW+1yNZ6d+4anMB5rB31WoxbOuN6bjI5Z1nbMpAcus/47p11w9bJaK3
2DVyG79cGPBtpQ3etEYSIXJgqsbnCeVcpMu5zPpdAWfGG5x8Ekj/De7dl8dKf6yqxQb1dhci5/nS
gh9pdg0+LobAnB0zkq6769+20SzGZA+4KPcN9yq+Sz1jF6kdkeatU/Dfk56JIrL2L23slnqW9VZl
/jBIgA17hu70VCnh8HISqzaigUMvz+2mvR+kykzRIZN8d91NBeSyPBCmozV8WFiDAGUu5HxaDsIF
+Mflu1DsdhhKNW3BlcRfTsW7MSoeXaAu67BoRsAyP6n5iNLW+a7ck44bl5hsbckL2UCjJtTf392q
vtVP/nVevbWIdAXa3aRb6RS9MgtvWyaSJ7hHvtVyqG7A21B4meBgMvfcqTrNoEgokPIi3OCPUCUh
cS2ZKLc2TVW1y+zYSsKZ7DN5uXJSL0tB29dvTp7xrdHWEa8JFE/DvFNO6D/vUWchnzkur9Na4EjH
A0PafdEhl9hVl8SU+uIa3DxIqToPf8y+LCea13BrXT1k4CmhpjYKBoIxJtKmc0aATqskFYTOc3JR
mf/dBrpwFlJUr/ZU7gVIWLl0wJkaU43DYFLTA2ogXWJEyBDnoM1sVW17yM2yoP3wX0lTmRZRNV1/
74jVzeOMXz2H2yVOFLijXDR49Je9P93F11myZK0ujiagJ0vLLrZ8djeyK3pD+i74aRwKw2BXqf7j
gye58hv4W9D2ReksV5FhdmlHvinVx4GNUyRdN9lzjjj+KkChvn16jqGlNNmpgC2pU/SZf7SJMqTA
6zIE7K2N0g9Vs0TRey+COJjT4c7dgtQIWSPguYGfatVYfXy4o1NOzSQv+Ebb5F6AHW+j9k9pbnIc
Yf++x+mBw1VQpNn4HD/OXppOa6wA1kwQcdzm9i46GvihqQV302Ecx7EWDj51/LumVbNFd+4xFGiW
5xOgb3QxGpM2gp0AYA6WuVQ54j2/8XjQ5wVWgJiccIU5MWCim09Jt+t0v+a7AL79HFv5LnJVBOcr
WRd/C86y8H9+6wY9j+EtOV/Tzq1twhfYecuT+vekB92KeYip42hfOCQ0vrCpyCndARQThl4wL5If
J/31KD1YytAbH69yz3CIRfBTLQGNDbFGbmcWxLSvQXkFUUkssvUWfs7/GFIXPVUoMZAUqwnGxaNP
cOAyYalKPGsPbYUVSQ6xVCd30d+vgivJ4LmTusS8ktqgxeBoLk/wzcnxUKvOuv17IfYRZo+p6Yd6
Vciz4sDhK8ogEea5cAEw8bZd2WrE137IEbRgRS7aBas1ldnCWKG+oNwgudo/TnG9Flf5tedinlgs
PMDyPvC9jxFoFOIbQYfy9xgywmwoaUxfB+9jAdk1g0tCkQmNYoATQ2K8HvHDXnOVY+CRmD7vaohN
FekI1+fl3tvLdlKMQ+UTsoDpTkJXvQaVRGkltRiJ1LGqDWmJhf5ZZijJxxvIJ4V9MuGSsBtmwQWQ
i5jKGYhBI5/J/Du+VXHKXPSkCjwgqj6Q+8/w4QGc+GjTLsRzXUk3aEilHTk224TWgcsgbg8deQ96
VD6V+/K275u0A11lkhLrkhi7qB3XcckAeXmi4PQDRPZTkdmjU+Z8/32MV170oNV+w2Eyu1/RJMcv
9o3VfhjrKO+YNn30Mqyf+JwaY9n4j0PjC4g3TmkMZe8KUiXXFOgjhaKjc9YoHPc5gqzIvUqGeBB4
fclu/0soJBO5MBvqpuiMjaw9Q2wAhTRgnTZQbk/IteqNOR41eG5c6HMnXJeNsG3VhLba/0cGQdJ5
x5WzNQqQTLOckp7Jbac376oe/HlQtQN5Iuaot38JVPtxlGxGt/UOSPXhBwnwWogOW5r2FgYqs7NQ
9k8jdZDPX/YwljsIPqxj1YBtwupHMHLi3rI1FusfV3y33zzH+mG+IDUc55BZB3g4xtOnml4FGaql
U+mazlmDrsDiyRZRnplqWKuPWKJQGZ8yqxumW1b4DB76SasZ9VZ2QXGxTvC8R2C824sO3Jzta3T7
ocQ4USdK85dGJHcMw0jHF7ZaohNFhXZFy+5KBGxhurSiW0RLXpKIh57xq9ATO9URSTmauHhBqCoJ
pYU2ms9pJ1RT5a6ZPWHe7Frti2+P3YsCYR2bFUW8kdsDZuDZWb5hjs/kai89+Qqzjyf0ODwSHhnH
/PS7KfEftWYYV6FUD9EE77talD1jhPDg1jK7Ii21Nnt/1GOxTlZuPquGiWwiB73fJxxWcuMr876y
ucnAaS+2O2fOCcQk2FMV7LGuPczzrWnq7qU8nPbMbVoQ6OFqBXHm5tTaLNNAOgwPny0k2Ily2u88
eK+D2/RZi9HIVCCSrWm77KPudkYyJXSbRObNrHwLOjsTSAsJfr65dqBWMElIzUQLjzpqXGMWikXg
qFFw6qwpNLYamvJopmGFEHrymksmqFTzzRRItdfRvNABpw2Lrs45vb267ER08zjbZDFlyfmSonbp
oHMZGvzzlIkDRqnMk4g/tvEZZAjyT1IzUCuKr/s1xbvqUJeY2r5QsGmt333uNGunakTJ1tLwwX6C
/ZdbfXGDq/xYhuxbsQUmz41yYzmanlzHnXN1GYW2RjjSaXQC3T52HyXTYobgVqo7JFjUhR6T7Mji
DC9rNKBNJbN7acq5ydcztBbsPgASFbzbZW8GqL3d/SbFJUJ2wNp7j0flyr2EZnh+0Naw5Ppwbwc2
IwjtKvgY3V06wp2XNQL90IqwkBnF92apbkKTEKujLRCZHGqaQAaGn4cgQwYC1VNqTGgZO67u/xLl
XR35Z2n1R3ATbaZTmmEVDyb0SJUMDX42sfNRGPg1b9dR182o5S7QNXCD2Q03aw+ChzLHLbIr/OIT
A5+Bjt8UNNkhb8MgnImuzlrYy2HLOBEe9hYgs9tfrSDMokwRYoVVZWZ8x4XkHeg44zirD4NCKdh4
pP0iFvmDBzeOKW6Hm7SXqZg8FXhCYViTDtYCLbLJlh7W6YbrtRM45BoNTSPz15yUB5qSxl9MP48p
+zfmmERLvvY5XPakmibXLLVxtuzEGDx/TKEKo5HdZRarYbQDdnGn/jN8EekHb+vNvvBF+enHsjyO
YDTm74QsHajV84i/n8EeaT7GC/P9E3cy7fTOaOVftubbX+WkIgVlJOPfZVap1dkAZQvOZkK6nI3t
hCetLRfGAc4QV6wsLJERrz09QWn9bAajciIemZftAWcMGCOS10xpYGllKLUfmLuyTFwi/GZ1Yu3j
tCL/VPqoAEwbJdH0TAoCFHbWU4xvbk9Ug1IXuOKyR8icafQrF/D/bqihDo/tzSjNWso/mUpmwcEM
ovkBwV84UMnOGie+ED9zO7IgqaMsieDDMd6Gc3IQ8laPT0vSD6yzs04ZTwy3LSrjfZW+3v+B1rTQ
Kb2KyHw9TRyIWMmB2rNct86tl6CF7+FRwUw8iyKsCDei/VtDnrBeWryhgb1SKNHnxhVSazjw/vTK
xvfPfeB4JU6XxS2gUhlvQpfSvb2yg1Umrl+drpbp8Jaa2aGgixAYLXclsyKmZh1Ou4F/EZIzzPx+
eYCdyWRczTzKbpnEqR+oq5hchFD1RK5NCPssGdYpSwviebmkwBpy9eNDy/1CFzOr8MBiOOpkOEKm
vikTZ7JSCDdsKtCqNCAFVxH60JYlQrksihK+P+CD3mUgpgvuITlhDqYo3HzZHl0o2pGdhsyB1Z8F
pZb7N+0padljIiMc4ilOwLvx/OYEyNsdPBuUky+uei3KV9n3IefxGx5udkHfnuvFU2IW+2nV72AD
CAejJQdtTOq8Ma3eGbet/BXbQcqooMm6c/+L+gtGY9fDOPtaGeMvHrRROL3ZzSFI8v6DVXjFHNNF
kvYr5qbbeZ+kU4GfX8YNNNuhrWA2LDobcwHZgy/2vHrbHNsiFH1Q7GA3ZOwdCsmEdVxDaJxVNmtc
wf7J1lrAhFKGNiruzvOYjrYTyUFdg/tE6iJjtjsuT9PX/9GjNl/PIpLcvMwn2ruE3pinLX1iQVvH
N1TN4OnxGTHKchpBpb+mkmfugU8V3SYMd87+PFCA/lHw5G7qDHD/LwkWF7diAbNOwxD1pQaxdJBM
ol/7+02Xxyno8yFvlB/v9GjbT2EH4gBSdVmBU1xuF/y3V9QTWwWtLHs66jrDnt+0XXnm//mfTX52
DGi6pGHvhGsObzskEQlzstF+6CL3gjQ1r+AVBhPZ1dZaMTls+6bjhDiCMx5ZYxlgLJCEm1zjZ0Ex
b97yn+Xj/YoRn1g2E3lXj2y2EFWgW8XEyLp65TMlZwj/3/riTR3fd9949I4hInsC9HLGyurXKVaq
7FxSE/+exPohkURISqtzC6oFpK2jOMb7tgZLUt/4DugfO5FyDg2KoBK7VsrZ8+QlQcHyQkmuZmMm
uCALxUovHVXSU1ukrjwmgBrHHdCeV98i/WNVJQG2vwkIaNqrSpOb+kizAmOz79KApebjX/da4y9Y
Rte7Ba1jjHLP0Hn3vaSCeIZlVffedB2d6GkLN8a0S7Jd6Bv0hvmtdJFSvvSoTvVy1Bc1vzjAH0xi
oK2eR/KFn6gNZ6GqmW+O5ofZCFoYlHs7VL/xJSFWq7JPTInG2MS9vLvX7bJH6ZHda0DZOg1ane5q
31GGqD/MAk7aUuJAmF4uVs7pKGpKsBzWvqPdmApqwgbsljjxy/aedi7DhXETTCylFcW8R9nYDnPm
Pd0l1RRDWSAcC5nnnV+6vDJDKJyIqKeNmMyVNLclpsgoIDF+1KvXXZObsz5U58lAudQgEPtFHKg7
vF6k8eX1+D8nipF0B7vgdwLt8K0c6PvG3JsN7GL2hX4yJLfw+3mqpgLZXjhTgj6IkRSlZpRoTtsb
31Xvdih/smlRITxIJUkS9NKZYHRvWTa0WHSQqrPuXdmzSYflmC9479X2rDBIsg1Cec9s/Z/pwXDf
xry2KVuTwn/5V8CPDL4cGxbqZIQL+ydNYfZ47DZqdWyDj4g/W5c6wmeqM3yato9wVYD1fENIXJqJ
54BTMkS1uwDtURtqCkUbvpIaqSwbIGLJPBcWFKOpcXmAXq+FpCMfSm3iNiKk22tgcJjRzDTPqfFp
GQ2+jqk98cybqZi+oupP8cFfqHDvsX5Bxp3vOEGlgf1ZgyKho0EpGtnpy6kUReV36lxZCmZk5wEJ
NNnOv74hEp9GmAt1819gvaHWFyMeBKyVOocaEt0Z8tWn5D+Lv7Sl1MUjEweGdFKGln8QwU30lWOe
TapVArTXU158zP/0cfNK4GMbNcmQT9LRuD6qv/VYM7oyx7pvuzsE/H47YZEFotMZd/6XZk5tWBo4
BgkLOTkrw8KUpZDqCPgay38rs71c+wbAmxilALJXhXSu1MgxwEfcHe+DhGlm4dspbvs02CK/ZRci
d/L/X5JnVLOceqYzmSg9H/T2n6mK+HYMLTjxx7ddy8h2KOq5TWDVdHkxyw0BiDXolBF7ZFK5ql8V
lcafmSBz3Qz/94w9Usax8lshTHVIFG/pj68JjILL9z1B0jzaCynPGL64eP1shtudN77m+xm5YKCb
jW7yVgEsi/Ic9REJarqc5VHdEb7mb1eI3Vr5qvxpqdcTAdgYlJ634jgiyzD2mE78g4ZxWorRSRnl
JftrqNhfgCiKju0JCh+3LpwNOdmi2EVGTgtBC6xeTmyzbiSysrPPJhR+inuLfGwp9vTO+BDv0SrS
9nTR6oxGVYGEfrgdCUXh4Pyum2RnZkE5eKPVrD722nhRBYnfYgeoTIbf3FO2xKyEWxQKKVQv3Hiq
uUSpstjk1tkLb05gdEj9bHG+FOLOtoQN2FFCXoNHzIUrrbhcJ49skTxOv1/d12i7CWWxPMPnCgXT
7hlJka3EdfzVcVOsD9Av5UtRAXqLolTP1U4vd16eQUSGm8iFmtB093u+FP8VCEMlzTF2Z8gFalyh
awCqYPPmGM9vN56+BnIwohZae93xUsa4u0iei4Q0gd+2rZ+niZgTDBjBsJYEeELvQn72Qqywr49r
pFlvyhqzg4d1/O1sOjAYiGayqr3qvFzDw1FW0sHs9SRoPuX0iqBZ1aNxfAFnLvNicOCVu7FaWC3/
BBxyEa+b53IA4NgCzA93+PGtjSQ91kn/gXF9XuycBwJErpmar3MFzoOE1PXf/CJVAjJfGH0Q7HEf
ctDinU3k92ZNHXx89JAMZqiMbKY+7242/BvcY0tFS8s6DI/OYaOy/j3O3oapRCIzLosvrvOOzgUd
2AP2Xm5//asiN1Z5C5GF24i3aGQez8H4UctvHK8yBuhUQ36ffp7+yHE9ZsiBmZlGIyeT+50tItkZ
xLNqNmgEXgLSF2BXLOZ7sBILtftEygzWxXAD/O5FyUpSqBkWzg9mtnM0Q4+Pq0Fk2MYcGNyBVe7i
z/7CdVbb24zujxJt8UIipPVoMCwsllJXJZX/Hr5VkUUkO8B1QJevPp1Xb9DPrIyPkFFTdUK7at4N
TUXLaupOAhcGyA6CGDhKF7q9B0z0+fzGuPM+gnYNpJqbA6ZoitCpnKtaqdiKe7HqXVWc+uyFOiUE
B639oIsUv8Kf/Ta7kSwRRwzlXuroYR57KVnzZ8Vpiuh1FNL3HAszS+ZKX6Z1hjMkrC2NUQl79lKi
jAGQe2cUB0w9Rjmapm7It+EoVYz8tQliod9l3tO4KDKqoZF+LBLra5rDYUJCt6EYHolxMu7ZYocD
K39leu4vdlyVi9I9aO5z98tf1QuvZilcLL4Fc+E95yUWYr/z38DS1dFC5Hj5+KV9fReBfj011pt3
JZbEOfX0rOfgMQKOerrF7ijGAgNE4ITeJAy5RjLxH0uvI4pv+osnp6pZFOkLL6gqVyszS1Hxbwwr
ltKylWPD9Gem++H+rIEtA1E8rysF9fFH191FBteym6yaQ/CiJjExF0KiLxU10bbB0FGm7VVk5vHV
I+pdkV/wGkunSJl0VIGVILMckOyJ5C5+MHTa+/Z/hjqRBcN/pFBNRZ+UEMHlCCZ6FmhnsoV9Jrn8
wwINLGPXI1NPVLluB1TIjgsqmgz8ClRS4fMeQAG8B8CALP0Zl5UmFQ0QzGQxLxNTDQN/hAXBw1JM
acrmVdH2WyDzsiN/uAXuYycL4e7BtQxu5KrslULUQiib3VcwCn3FaBQV1a+y/ZgAGLu1jxjXRFdA
h+ZsWq7lmTLlE66xgUDKfvyYjHiiuQJO7MpM+Mipf+2vpQk2piROOd4qxmO2JdM7M06kYGooAyV+
Fxyf+pHGCNsYWNx6nL+si44p7mWCrRdBrVk3FgnWfON0XhwEpbpe9Uci2GMeHuQdGqrgDpjduQkf
UqiQnbmFPo8t3wKiIyfWcJovoeLLLzQo4x9yuiACf8rVxO/UtaqAc85F1GyQnlFlK57rKcksgabH
aaUuXS/0bJYJShe2m5i2c/DKnPXevy47KjV5B7d7uJGXdGrgbbjR+kywZ2rITwauTpu112VXcDkI
mJz2Tp/DfG5DEKnqi+M1/jqU67IGTfN31dYJsGzJKDvUwr+zJrdshK+Ama8Ye+yT5kJ0V7Q/v1VI
vpYbGM1EyYv9jfBFQYPZ2Rqy2nxlxHHqaLgtBLcJu0ggqEA2jisBbWY+wM8ipn/dDYRLnIlXxtar
MtfX048NIN6m2nSb2wgg3A2hTT9A0fc8zO1VCtmX0sqcVcAT1auH1myS0/GEHc4q5TbWYhIqBWoA
SYOVT649pPVgw+UBbUvtwPPa2hPqGdIX1MU5Tw1Rhho4i4oUow5MGtuc9izcyPzrBCTNaGbar2Eb
yshTpUzV6yAJS0cajEolJC5GjczCrJxOl/db8fYiDsPzr+Gphbt79WFjUQkvbsBMpkqUXSXiDm/C
F069vLi8ld5cOTJFqzKhXUO0A6emeSkBgqlTavGqcPfKABab2fX7YoTroWzIcMm0uco4p3sAoVJN
W6fycWGSSVm7ylCYSpRlr/5NHRsV6ug79lbGAi20kPl6bKeqNlXHptf34IA169DyJ7R1/ktEIpF6
yVtCcrpTl1mL2YLWpx8eqPFg1urbQsRQohtDXBgRdoFi9vuiZGzVdYo0AoWVnLW1MDyTFsDT9F65
XBn24GpyJI1lNwdskhvFOjHaeSAOiq+pR92dWThsOJL8JDycyy5QsknYWrQYCLx/u80x8sPVkiMQ
egmTIjqwOOnuJQCXSkOrY9HGVWbbLt5INQRVXJUywJo9vAub2qtQrVhmAqoTaSaodAERrzsMjjmD
UbsCMItZyQ8NLGt0VH8i93Cp4s7IRxBepMlKcmmsyTQa/yoUzxQvEWA6tlCxjrquiExAmyckTkqw
VVQoNoE8VY2PvNJiQNW45iLkTY/c+zS431kTaKQTJWpyjfUFnDImp8eYhHMD5Nq+ryG2sYG1p7z0
mwkyb0DDGYa3ce+18GtUx5ynQJutaPF6yg8TE7+qYi/D6ZJ6NeH4qCN51adqbeyk1GqA35PhzEyE
hl+vnJVm5kswbIvUM9+39/ZNEf0mTcm6PODA2C42IrvEALDnbLh7PxkqG4YKyE8MOfCxWk7lFrbw
T9Pvnv3IieyqEvUn/Uc8gWhso6qQntUz/6IE0udhFt055wG2pJWwn6yzd+ztkc0cnSHO9ldiXf0b
sKlSu8t0RUY6XwQVpKCb2PXGx99NBWttssDegRF9ZoaAPkO50/rTFRPRS05YiiaiEwI9aLvm5y0K
s8GatObp6kLg80OuZHC4nfNw09jOIqFdGvAEXPEH0t8i8zC0cd0Rje6QUb8DdrTjDTfqJTueWNz9
3W/ZObsEU5gawscBjZJK1SOwQbshDScSuh2wmUBa57EJXUYHwN9A9NP8O+xj/Zsud5IjlrpmtQVw
6FEe4ggFaNa9ZkGwSejPWQfsu0RMMB/VZ2LN4ROItgr5vsPpKaplnVz3JdZCvIdJ6a674i03G3Gd
UsCU3nZaZHUPtg7n7DRJ6m0zZ9Z5p7yU/MFURfNpD1Ph74ljRpsNOc5fBq900mDkIdEZ1X03ybJX
EV5lX/igOruPPb3q3BfNpcFsMAyGi9oBEzVGerybmJZ0zyMict1lW9l31it4r754L6I47rKNdT4L
ZgSzPTe/AEyUPxtYgcGX9ML5B84Jxg9CGYuNlCrV/bTL3C0iIs6sq3taZezC1oO7KOmT4tGt0C0K
INcPgod9Jh+7xAAIfuWZ+D+mUBk+WUAPbQA9XcDbcGsVDA6vXP6sEtj51WOYs9lxx7lWvyOQ9PVe
dyVE+ZQ/jqOkMuo0Gqa3W5VbPFUdngaXeLdWca4G9C61lWMdCekXPve/3PZMeoXezZeaD5iujPgq
YxEO8ZNpoDTztG35IgMPT/WV0wxODae7KjlA6hU8RAINw/gB8ZpzZTgMYVgSJtFQCQ0c5PthoCDE
4gwisgsISrOmjWr4v2hayt/Y4hfxSeTjdgmbLAxpGsbr/hxyXVlK0WwcLAKA/zG2b6pUvVfLcaac
KtP9TItEA0vywvnraLYsv6rG39bvAdz7ykvpXTrWlJoEUcK8WPBRY6fvti8EdtvpDh714T9nGSed
/9JZy7HDp1dV2XFxeLioUkeJXvQOWvQnyDGCQ9O0xDZbEjvc1N9+cytUx9mljvMkZuGJo2fskS7D
M2LZAebsaVEynUbnXkxzxSumTfZRFMGzGv0W6LWbmrBhgjdb3HOeOsotwi281c/BFDxd9egVzDWd
ceJu1wRwUu/jPWWHD7pwHXnGE+wGtr9f9+RfAMjGg5RV4345QPlXduATQeK02ktQTb/9ydevuJZS
4NTkribRBXz9naeijC4KPzqdyDWrpJSMiCabiOqCmg+i2f11nw7G+fd+s/tneDUAJ33xWLpqJIlG
hH0IU3O6Kuz07QBBgqMXwdAezPt/ftoUUsWdSh3qhbOknVhMM22A/Goa3UTfzx2d2dy3vYzDNhaP
cquYNabGwPbv7yrJ3z548rIqhYNhBaMnCZ8JqTx0pPEEpu+Z/PcmIErnS979ei060aaELPznj4sm
r8AyQ0LCYklt0kaxuSacqdKoJkvpJavsPTZYRUGJAjtN1GyWTcYEyZZT4eFdOGJhq3Pf0K3UDIHU
bzyOMPylseicvymgY1oGcsN49598hmeXHQ1YUJUw6W7c67UKYA14yRQOQ9Yh9wI/xijpscOtehqx
kDXV+7BqcgGw/pOgDERZ+0ULbPNMbLUCFl0IQN5YHwkw73g83ODGmGBbE7rR/xPZIw2hStZUWFwe
lsqyl6eAsFuP6r/BkRWiThUkK6Kt/rpGQGCy8+TzAywAUxKVofsKNOXr0JcHFoC597XoqwDQCNb+
Cxkzwp2CKWqi6vYPzTwRSTxSTtokl1vxUGD4k6+0i1lPZ0cFVXSqsG2tZJu65vJ6I0nwvwDwYznO
8DpIYpl8gZNBFzv8EtKcjaJUau3KAJ2TZnEXXcxhFUNzRCRNzS1Cc7TM+8ASFvgTVwqs5DVKPSyA
i44s1oJAZ3kGJxqo0IR1SeCzPEFqz2z5FOvywjxB0ikBqkXIDjnj07kgoQJcp4qTfty6apHhLYMt
iC6ReVt1piCn1LuI0wn/HiqQwAe05CnWWR9gXU/wmax/cM1htmDtaNUix8sKtNxAJQSQ+dN6LXZl
wbXhH5pZwkST1Y4u3YrWAKnqCTe7TfP1qJblDw1MNZT0mh4Z21tsMMyTkkhw+93Zrh+vKuXVkPs8
50USOOr/vhEMSDt94jGTrV24gNKzW7/YbuxoX3gKAv/l6+1DhXIImNvvkIN098Lm0jjhfGXX6cpY
F6tf4umQjiQYi+XbLw4cgZ6WaQCJshv0nXgy55+rSjQh3bEeFjgH02po6PMWKjjzKmpfiszvP0nD
VfjAdl+OQahWS5YkGWFoTBEEmj4USyxOnDh9QM/rZcn5xSMEhMXGPKipw3odv0jQ6fMzPN7gieiV
/uGQBOupzKujN21GobiVzWxhSg8tR2t6egMbFxkEAkysfUKmJbluyEmjawygWECMKA45/r5KWo8u
Q40GRm634MKuifr3cJnQdVNd5MDfTNggi2rTMiX6aLNz1sNZUb9uXEx+PAoWBTDL1XTYHH7MG4xw
bhoNqWR0KZVBLErfxC0KMnP9MSv8lnMxJCwTNalgOwIH9Nzmlk9usqiwJvxXdYyZnOudpj6x3jua
eO0vFBair1Bcz6hrD/v10lq63WfxCjjw2QpR2WkNvfV5FH4Ksbo71bxU4gqSPUKByhaOCzfa5V/U
5jF6V62RLQpn/QTS5hLSpr4H67uk/8melHUdJH30po60KEWaxQEYTU5tMjgXyvJ8GaHTr6VaPx3T
xKJ8oCa6hfIsE8GLQZw6BAVayQi9fhtG2BGi0Ss3wn1/7Lydx43BWis1Z0QcznjSvu/6HHjyxBjP
NowmNTB0jPvi/pbuK8gmsvJ2rZ9hC3SWW71iG2GdnFNYTWdk4zLtYu2Co+TBkIANRyXyBbveeQAU
3mAy/wGOuxABtXwmusc2WmRZaiyVVZslTzsg83ZZkO7Cp8uBfKazqF4IcIuESadUs59zQ+ZUWk8D
7NThlj23McwNbcnqmoZAEqD5OUlaMtorckr5jieKRUAsBKSwMG+olrs264JGSyviu0F9B++je/Nj
QrrEw+9WOVk+fwr2TI8N9PgXGj4rPUyj7rqoEOc6oCZGFx5lOSHk+MEIc+UWy5m+8TKP5xrNE2q7
No3NySw4x/bA6wP3obboYmz7oMd2PV9/k96AKGn2djA/7sOEduOoayV1yxz9ZmGsI8WUtUUZ45qT
KWCrqy28SSXX0qUxDsvxQVjAu0TGnx3mZVYkDuVuG7njAlOJ4egEWSaoOZFdMOTavkMLZR1cln02
RZWaBxHZuxCej+1JSJFvTmt50ZXE5KHJG/HI9L8upuEq1mijHQlSU7q9LH++JMJuCxrWgF2XAadv
ZeosiLMVWWlGtz8huFuqErRM5f5Cs6EmLNkoRO9HJ8CeynWoCYRtTo1iIF0Do/VnpLPtKfQX4EoJ
OU4AhVVEqKvFFoW0jP2wdxPP9Wd08uI7+9RhEdZ68O9XzVae0UmTyI+WXUgUaBbkUQNnL+aC9ANo
TdJ1b86i4xjP28BWqbSxpik56ke8zWZrYAE1iu42d5I/txm/5ANQTGmelITnBPShjgLgyIdBd0ai
IuM1CmBRZGtJrqZncDsRvLy4cHQkJrKKCCWXUHGlYU2fmw3LozlwdCCO332DNJEcWhZhgDLbtpUu
elhAKedpcmFaFd+q0LrRWcOYXfDPkb4YQbsgReHcm7DOk9Zpcy067lL4G2HrMLxt/t/TG8U94/qw
3jgwUzcnfi3g/xphC1zruFQhnNTGv9HehNtnOBzR629bc1hPOOYFiQc6hrCvndTfwl088DWLLB/P
JgDneuSHByxievC0QcpGlSxP8KzkcDQUic25dCZ8N/coD3Hob1tgwpSW0TCTPRma0ANqyfj4XePj
BqCylQezTed1vfQGCkAw7NoxIucyCXJvnTeiis0A4uVYPbBWSzocHSsQnMmP702XxJx3dKleFuYp
2dyMrKMnyyxVba+TQQWPd7SWITqnok1Y8Cv2pDEc8xhve4wXB3PTL4FQsyjqOOhIogMbubpnFvMr
ad2q2PypWJHZRNKvqZ/ZOKJJCLdCA99sKjYV7ovkTDGiv5shYc74GYH83JJ1oLl2DPhx2MMCutC2
AzCZv8Akm/BGwxdN+QEa4WRaozKu4woEpYXrtl0SSOqzWZVtVRBqE1kmTqH/xaE8Pbvrr2IySWR7
YX796VmvtjEPEowro2+M36n7vVbXFbTAl4xGXrnDNu2Qq+oy/zP4wmGzbwUsXOhj7kxhMDzPMIun
n4KbsYIJDGfByPEj6glYIQjGWqYMURGP9fT39fJ6da5WsmabaP517JDYxSJwS3Hz/s4gCqIVj2q9
mGwIYXoZ/sDWOAzXYYKszaEZJXp8QNU6jTDpsChJrHlzWL5AAMF+fy+ZFADl+I6MbaSnU/dgPY8m
O0xT67UpF3ZrI8c9sVUvaafMpqTXwEnRBcz5kSJJ375D00DgmJ8lPu4P8zlpODwTR2iWGzjYk5Oe
Zz/fhLts9yGI5lVJ0A1He6vASM4CEwNm87QkGvfV52htlRwBJ5z6nqUdF5IBVIH+KgNQNBNVvhVy
Vt1EB9bXG9heOaYX8NYUyEukeXtPrSC1qkKB5NfDBtZtjF9fd7rSUIMXRY7rbWmoqIM0S8lEOZQu
EB8omirjd2LGf3F4tBqVBIUFVHQ9cZgziS09dvV+CjGMQfZg6LZtHhFnDcp3L0YpB+kJTUuRMfYK
J4kec3EBDDm20na/fwYNyaAaglFIhPez+WMVehiul5et9k3DPylOWOocEGLGjV16VOr25astz1e/
WqEZA/sCaW9Otn3nB6ZOQf2kcfZNKbIyXTAfI83o1Bxy8SmqUl4wFKAcWr+SC+gHW7rwMh8biq2z
LaknwwEzPkl7ngcizSP3lbdeWh78Pmh0WG5R5F1YxhHWqrexlnAYttXkfHNhGivsYIKY0uR4Bdjc
IafozV6n1sw4BAsNx2LSZMuor4OeAARaXb8suL4qDXPa5EG70jQvB0PucjRM3IkOurBfrA/ttAmT
G9mPR9qo4a+DaHhh+IMHy2KgjSo8WDMqQJQPNbnAIIsphPq+C3j7SAVfHjMRyhfINDdKM6OSURlW
czPZODHxxcuc3o7JA+M9PorSKugXur0zH51ttK9QVEyVnE1uBETlUjdp4wd6pm9f5PBGilNZb5v2
u1ozokKygn2EhTKzIbJJOEalvxjuJLFa2EVNB6EoY4nYDZm7KPjQaa/WSnyy8fWnxYQUiip5inGM
l+xqkmW2q0doVX9QdyCRCAhOIIu8b8cUpYuVrcRISQxYAiPnh5tBaRz1oozgxQdi9673+1xzOVpN
5d0hJ/QgMyAGtd+gXylsx9vXVHdCDi76EHoa4st4pMi6X9+BpBRitDC3FEstA5+HmzUdKC7XniNy
3vIb7Ne1RxyOSFSch7NBXYow8flbjsOFqWh13iPvskZFDw3ui0OZZlLvGCVNQAIA7tVgbIdpe/FW
tcu5Vs281q70yUPQe1hRZfu3Ymkw5vSwm61JSIMkW6DHJ2Ouhl4ftJNhRU1Dqz9RNHjWVRbUvhj9
0CK16FzKLCkaaAuTo/WWf4LOdWOycgqXQNi+/Y0C+d2pAaz0398Rzi8ZlcGYBgk9XY1Y88R+2DDA
JA0JxxyqMDVXCBtjglZLg4rxpoFx/6pmtcRro1U+h5EkpIjxJ59gpFYio0TWPA008m0u2Ul3dA+P
WC+OW98CtCCzvEkYztfKFk9HNxo9G9W5q+CAnUkkFF9xSmnnmmWZQAA1W147vhA034L3PR9D3P9G
6UZTzXKF2lRXu5NSWjCusKyvOXIPpRe3O7pteXFWu8VPkY6HFRnNqB/ozX3U2nMupdv5EDIDstlG
pg1BJikzWVbtcvPygiSLYPcjWYKe4iKFhCOld+hfluDNuTCWorl5elZzMqbsDmy1DvQQDT/5rkjU
inTfYhLcTct+O2YIUIxz3HEeId72Fws9x6JmvQwuQFrG3IP9p5DFHzHE1mAJt+fu89BGqoLSUwRi
kST4n8bm89/JHI2ekYKQQB7ga0u5StY7osIL3XCaT1qtXFE07Zzu+v5eBX1P7OV8K2OLHjwSi2Uy
7JM0ZxEeMspDobNh3Ysm4VoZu3TiAg7SfWP1pb6fhpbiC3L3cw1+bO9nz/Y3xbYfpcXj9uFjOFOQ
zH1t05NfjUN1k6AOPd/Rq0rc98y+V05b/Uc4u5d6p9kPg22aMLHAS1g2zN3dORYjStCE/93M3en9
6iHuulow2m80Np+25mCrNs0ypBlfnE0BdFMXWFrT+S1cNqbho3aP8rpNQpIvlS/5rcgJeXvXkT6k
bQXvqy8Z+C12v/nLFpLGTBHZ+8PkIe7c+RerIGzH3KQztx/VyXP+FHbfWWZR/sYyzehe058lr6s+
MBRZ+EpwktVBvcAV7bIio9I8YKO8VpwbNXke0W07d6Oce/xY+JJfFtk9L7Ok6YS9H95P8L5ll7OK
XN8yAZ/kZO/jlYR6G35kW4JdAHiicYvUgM70qqTkVk6PdhVfs5gCRmJNhAczjk8cKBmlvvI5qXFD
FlJiBdB0qfR5VH+G8XeyAmPYH43h+ItVVeZJyQZJfGvUiW5g/NNARECG4p3nbV1FiZrEJXm1j43q
Yv2WxZd5en+4GjhLz7oH1VDmvYwghEQU9fiZzTGfcqvBp4SxW6bDYP0u6vb9hUMWvwBlXEPctjcG
KYX68M7H2BcX4pGnwA24wkWssRrj52aJ0eQBXop3yzV296SwTrLotiUUu0zolU2Xi0tGT+7oumjg
5rDcGPRkfo3KTDRXgzczzBhqBY6Hmd2FTjq+87TMKvcsBFjiZrT3zVwoVExV+DtZFtXSvVHVoj4L
MSOQTU1CoBNfHRsiCR0Glu9XB5BP62RQaxT1Bm1pEqW1OXsrnmICbBP466y2ggj3JKQ56xMENdN6
AYV6yDm0z9aD6ZpdUMIwo9Y2m435tP5CzWgcxkUJHjHaeS4ddCFpRSS6SQO0px3YTiINFG+ezqvM
EVKMcHomPTx8xPZiRpotsKDBW6ihWnCrJkhNwaJv9bZWmmHg0wT+ABkLKpUDdJgCc44srp105zCG
J4zWy8g80PAO1xF5icM7PkZHu0pBqf6rxopFr1XXgeUn7K1eXfI9Q93Yat1jmaZSgEtzey4S4Isw
G0ZaxpVwdOpDqEJVAm33a7MV2IFWmcfLBK9wpSvBTvUqdt2vjX8bQeXbOg4jQ3mo+3tqtaH1NWxl
ZPT7NZ6y/31rWR23coLqxbAht33nbfek+lycBqiAYgbGdMiCBL5k7t5SBPY+sZTtYTLYbkM5tufv
uXzJWEegC/n4Y/tl/wIRp0tWaMbZVeSbBPzclmqv8gfSohigjTSXApU9+TVgsaY2RCkNAoH+8LA7
rrD9wJpWoRJV0zj6lkqBxRvQhoieSbfZXoYD6ikaHUzye75+h1U534fhwLlD+3Uu+wOme6C27mYE
/b/+RNa7bObjqGgLO7gltCyXFcg/wqBify3A8oy5GX3BRLHbmHU8lDxTiuWkzzR/eTGWjj77j9ID
jC6vZLQvlMvXUgKIC81qcxiygUvYiJDSIojwXBqyTcaEUgvIeER+GbtXI3T7p7cdOWb5ii54OGzp
1b97F9nfitua+T8kG/9Tnx6D6Fu0WZ9G5kzcN03+9hA1LlExmkePSIGASUdJk2uDFF8HwQAwpfik
tnm0hBGVGYbqgp/K18Rjq3z/vjwYLhJU/COqhIMJQa6Pwf9xmL0LHzl1XzzdRZbfP+shLaZ8ZHad
UPNzp8TGFTZ1gYNLexy0eGbogXLsZWN77ezpp3/qKW6YrMhb6yGFD9fnx+Iap92I8uv9ErsAVZ8t
Qkn6/+bNC2lohCMR5NAsprgmjWDD8tIc7F6kHBcmqFEyZdKH5OHFZz7DNkXlpgoI/5vVVb/dPlwv
hIPbPP9R8lMbfKdSR1GI5I4Ie1EGpAW+EETq971E/7uR7el6jGijqhWfF8AD3ZApCLv8x4DIhSmq
g9Q8ItHqX4otBnFN5UAFF9DNw45fAmPvgFA1jBrHDf6/KrIDvk/L5KJoBNnSEC1JEGOGCpsRZGYS
WGmt6ZSH0jGocaMyLLVQEw1gDyiYUFdXTePKdX2l5EwQtMYHqabT73Zvntg01ubvKqtcZJxMp+Kz
4C/I8kbZ9JuQ0Mo/hekXYy8kTlgwFb39yEnfvrz9sMdZSrYXWBCdA8A3G8lNbHlwNDiQ06JNwSxb
7j+5UoTSZhY8pJPRz8qeAOrnzcIi6JMrPuzXHrLSbHF1WtmvaBu6nBVuJf5Cs6FTOI/38oDuwe1B
qqwfSFcLf5u5OHlrvHlJq/VQZzjrsbKsA5rYJHVgwOenSCRrPMVt0p1mRSR8ySUAlhlAh1OfW5pL
UhoAYYbUb5C91WJhKEY8JzeYqMIqmaWZnXiS7q+/yt+QhnlXytujXGCMmWy+jQwHc249V26sfMnh
hmNQaEd67mhWuyPTfsjf3QPu7sIn8J4cb72s3EzCozIY9JB9BM0cLbICB7tXoOenzBQxBDgrGzFt
/Nx+WqdG4Lolw9aG/10QcLKwkIt+J9p1xfW6oQzS8a4IeEwfws7LlwCwN2DKwMdtiAjClsnN45pd
Svd8LvSv87uhzUTUJ4TZFZqLDiSgFe/1B5tf0vVvnTtZWyZH0hQry9mP4W7oVqdXsZA8M/kP4tcc
dPr4U+9DxJEauklOiTlmZYng6isGox8IqUODKCrlPpOTqKoe1h0VmL3YbVt9EI2Qjzmpizps5MhC
WjRpAtjBLwcmHk6pgJRzQDFqJ5o+VXz5k9hshXzjzKQVIpikb/s7FqFfSaoQqzVvg9KlXPYZHEbI
ORRI9l8WR4aDjzsvb2misQh0mpiVJkklRHmkEcAkkASuK7X8kS5QbTQQSBrGDQn8eGydaQG2/aB6
ZvwN14RtXkWdEzUd0CGiTWaY7h3L9O0GHrNLbUXEJm0T62be+oErM1j8Yn3uGjjStBK54vi5l8IC
UnXrER+4V64EbQCNhNVyKEF4E5uTP0uwbmzgGY8BbYxg0iBtTJSHZKfRuYk4eNardKmuYJ29E9lr
MUMlp444sKz++BjO56MlTAi5wu8UmTHwSrHNKBEgoOcRihGjbR/eLylTezEI83WI32zJk0vIORb9
LbWpIv0Q2QSMfiKjn2KAF/W+4Yw+7HW3uOUQD781kuTDSiFQmn1WksKdLykgn6YBzEquiSEJJOCe
/Yrk7C2a1EaybYwgPWpivFWfqmNRbfhxVSyzxZ7UfNgTWf4w8ZCCoJnaXdus4rQnG3wLiVeqeXtV
MwkuR1ZphyL0kl9bbVbnD2bpRzM1LWqWttCYLU+gVXaptezw48725jo87HzSt0AVs9R+7zVYL5ad
a0IgBwUnQbOCzyR+vLrKnJYHoWpVO8frwIj+1yEeJwlY/4V17tPFYi9aQ5GyFOxgb3ukQ1/ypgj5
So9AhXWYVM06ABZ2GnxZhNz2kEi05z0jHdHOw7yWerE3+DIYd1AUcs++d+ShdPWbF+8R7mt1lzVX
KhqUDgzxtg7UGu0WE4cNQzqkcoUxtZX0uw9EaDZ8jWCnL+4H2sy5oo+fG5QtMvoV6+MAGU/fDkaR
uxeOtN/eSCpnzLb/E5iw4exudqTPVaP8Kp1fpRveOiuEo/b56DGiN3b3SrQUeWj4+HI4HAhmUCP+
ve8KESu49pcAUf/olCHA6v6BrUJ5b+dgxCf2CbRmM7wZROIivyeDPznM9Krl3ZGhoxzUezG+8RQy
A/tUVDLMnfUWctIPH6XNqerYRYMaIqXFI+H+Ua0avOuJKC6epVaMU5F8F7PDgwMiWRHwkIXYdWBh
i3kDSQnwk2gl0CcE6bmhTFxSBHnWkb7uu0h2JeUoJ4CsjeYeN4UQ8wcv4QvedAN2sLkW0JYo5bBF
TYSY7xziaCWDBgfPzb9xtCKVVC1jR18ByqocllduK1gcOsfcysf8vghx/Zoz7s2oE1MMeIzDfG/6
Ipj12VaH14zyZejanQ/c7tQHKLnxRwoDUq/439BJiPNA6AoDzMvfrUTVqokZLys29iqqc6+Bajds
aeQWBjs5RQDQZNIdDsZBUwaTOeHg7TnDIxkLRdK7I+NE1SR8siQbsPlrQOf6Xhlc2Y56y+eo54nD
E5Xy9P22DegOSQOJAAio30eySPK//VAAD/qyKco235ZR0BurGMBPbROJh2TbLRQB1kb71bNX6L8x
L4+8Flt5ymn0qvryWUoXXp51UQ2nLLtuf/+0uZ8Rte0/b1vNX6uEkIC0VTxuywIre1gIMOPcX0WU
RU1qJQx+VhWZPB3XO5ORL+9yvwQB3TZ4XE8gCNhaPkwrvIWjoU3fn1w/1yRW5/quLLaOKHIaduOI
+xv3ykghArycZD/8xHQx8zEvbpQx4M+WxNqhF/Qggw19Y3o5hmyC4MpZaaQmRMDR5dprZCexyJ3K
UJGexCyjZEL57jVIfs7mWAfpC0HS6RN1jRF94/ORzag/YQMDE2TqDU12VJOLgE1SC2V/7EVJWu6P
OEzFpRImsf46qLCFQh+rKsCPSCsEg+w7saHHhjVE3+6cS+OrCr11SzQNFkELZ3jGLOUh1hBXcDWE
TTIUb9oC3VhNoFVuC5+5CRb9d0z10URaV95DAmYAKH4kdvuUjCiKnv4nQoKE71qYy1C3kejpp20t
Jx7iQnx3fnviZ2mE04jki3pKVltOZ5AyGUdClfVskNB3FnqLplKEHNAr1b8BUIWQO4DesMxHeLgO
v0mncoRFFN/gtXqYgaGGs12KECiezYVi5O8fuHWG0EgB9tO2Kv8tT7kDH8Lmsb0xaZwXsmXCOKhL
Gc7KRLlAXtWsZmwOI2TyQN9K8xvDSoI9LXa6nBjV/o9QTGYzYYm9JHp9mnYeCUa9X6zMB9vWvz8a
Q7UfEP5G8WhsuSOgJ+5w8VS4A9Glr4Z0IrQlP0/xTSnn3PJ2nCy4FxtbcZB3MdXnvx03Sj/k/bP1
1Nq7m4BcJEh+6FZ325W2eNwl912R4nPOfsLhoIV9SRg13NIbWJSGVMx6GHown8kXdXmsDtvE0Rpn
yEGg4Y+PDP2BK793U0588T62Pi7+qG88yhu7kDypsWwbbcTD+ymQ9C4V5IyfnP4Aab9yqm8wuAKX
HS47unZat/ci8988DofiCXI5a3yBsdUX6pz/GqY8MyiCmo+pMcVaHpNUup8dp+EzO+nZ1cT+TlSt
21+lviWlgkdaioEd8tKxwfgAF+HAKOlaQveep1IgD1HZe3F+TnwF6mXxb7XOWHvvlSIXOrLRFh0/
jLVB5bQVSkV5FhEDVLPvXpe+A+brfQ2zYC3rTtnr77axbaeQjMqwr/wc79fx9NQiOO54/nvTiHbf
J4Qx7bB6NxNXhZGHZZGaOCcSalRHZVh0njp+BJVrwGjWYEjEaiRLm9Gd+FnGBSd19XHOePpq94yT
nCj+ihGN0wiN+lkcm45ODI9NHO1mra49wiA3TwxhbW/ekudZf1Mpp7KBiI3YZXcRCMhfRkmOowBR
LDtkIi3DlezugOQKyVgkSL2CuAQ9ZBbak9hnRxhQpn/mVFI4LNlYt7n23ae5C37R3VMQLuvzn7Ry
EQ4a3r4W0ixDYUx3bvPaMbJTq8YAqiKHOjFdJvhfQfEcPEgaDal30nnTPNPXPbs/pX60h/Z9Am6j
J81OAFJDNWQE63o0xglR8zwVmBdiRePBDTdzyCjn0z1ydZXGK7L3kWuDXiezkO+661GCzyhcqQyV
4P6U1sr4CqZ5i6PsUmvuiYJfF88eqy73kkytg/xZY+HJRjaYIrimERqkRpg/2hU5rmsRaS/fUaPz
FBj1Sz3m5X6WSsYVKRSHjphyRfyoF6UhHWdN779LGXXM/o5spIzsAQ1Ii089ewLVI7kNod67MDTD
DCi4cDOP9aomdEZ9F4r/elT2t+8qk21qSm1RlS48j5olGqfa3x2KmCEYcboh5rdxkp4m1kr53iQn
L+LiehwrHgkbCIijiPivtNNhaJGQMIaAVwUvOBjbRXUY65o5QU4rdC0ufEgHp45/o37zNvt1VtAk
KcpyFpgNTVTqwvXcDnFMXEd+lV6NLYqWt8H0Wn2V+iDyFP+J0obUnYMHzgAK+soZz6gV04jOWhoc
04XOcz5JTBvmDFN4OP/PaCv1bkx8PZSJw11pgGIQ+rZNeq94/try1pR7YBBkVY2oT6JeZsXV95/X
pPZmvlh61yU94k7doI1f4pa3+eU2MskIJuq16pisjWLonLXbqm3WuLTlbZU6JvMuLEiQm7fo/iC6
MGkeAHp6xdJv3VKIZo6vJ1QVRdp6e590Qqdgoh6D80cFv5lzirn/s/kiJtPmBvBB1VyIp6sE9FIB
0wlLs0UbvSa8YIJ9gAajviMtmlkLfetTdoQBPtkT2JPvQy6kKTsFR/w+Sh7JnZUMvXX5MJAGYNu8
quIpEBOHHH+Hc/CO0y/QR30T5wAgDs6VhXnwlAmeXRxS37S9EI5gPzTXMjNZkV+CbkIR2OS34dDd
iIIiQCNzoUnnEtPN3+F1ygM0hhiAzbx8Lz+mPasIWCYfg1O+h/x7HiREktattsHRkANuTQwwKK/C
rnMBCtLkB0Xx1zbBJIKRJqfHzTiC5H310nglqicWrKSgivOVU5sLSpzMt3fSIyvd8TCfusa4b9zn
yhjGtuR58OHt6uEEb+fly9EdCg+3AHe4tlxOQC8fAClTvLsBXqInNKgQ1GyijTOKAGEO4aA73+s8
0cDQMDxvQE9j1szzZpdoMwX3cWuy8/bKq4U5+5FhiZCvMnczv6Fa/KnO9GI8HHkJGtp+5XLyUu/E
Ie9lMbgHY5peO3ho3VJHGES9FQSLwVJ/5zxrOkcQA1HL5yZFDiVfHUetVQY13AlTrHuOUgf7H4Vs
BSVm8q1aVPvyTTyosAvVqOFFLNJvwDBmR5c2eqyEKdcpAp6466E5p06G/a6t8riQL3u9lLtnD8zT
SNUyF4KHyRRWc3XJSVCepBERgU+Znbg6Mp7eAngWrtDfkT40vi1uzNvmlgIvp0oex0NKj4wKez+L
v1EJjvEKnThqCRs314B19W5LTWUBlsYbU573AfRdxTCMFf9O2loNONevrJiqaUIAqopfKE2yT9kY
RggW3CVUrMaNHC7ny9dyPgJdB/Of52xqUSRSHxcaqk7umhp7TkiLIbiEFvqbYwLSboWwwNt+d5jb
4ssXKw7mNbAgpzKaIf/ukbDF1F8dd6+AjOxoU7YcgEATy6QxaxWvGe7Zh9jODpn2W0A4FLdj5g8s
Mbia7yIt8snMsFHSGgL/jqtFVbh7cT+470G0Sj6/NCpndMBtMNVaMri0NXh1WqnyMyehD767Lfi1
f7OMelqC1c/JtiIxQRt9M4ksB4odkFAZqQnfXbEpkNStwtM2C/A0rbkX4xucibW/VW/LJ+41Ix3N
elWs31SaAKZ7ugka8YbQnJ5asIRhIsWjIwtko8V69LIWQn6ySLMLbFsFurFfKLPLkVDPCGOxnnyZ
4x98u9oUrYMQA97qVDl+3qfO/OWXitFDlEKLJB4AQheoZjEj8A1ehrmhUmOA4cnTP+qdw2/r0Lat
hddRGisBuoyTyA//Du6HW9zgCwJC9csgHWaSejzAeQHnnUTvpxE0mHmOIxC6eT1ButQt6bz8CXDM
9d4i4jljFVPBEAqyhZp6OJY7scow/tjH2BjsoqpWDAy1/GazpSmD+KV7q9uzWX/sagTQlDKMPV/+
hDRphmbLtC5Gjogq2Iu6oDIpAHoELHCAMekbrpOc3GHdoHiahOpC83wkUY5Te+NwOSmAwxw+bIs3
wi/Eqaf+XrUrmbIZqrqOSgf82U4iurkjT3+EDsmie0XexlZINEz6obsBvIHbuJAyNqCjZ9LWrUBP
ZeSoR9w3DkmY92oT7kmhxbFYLYhNTzIQWKiwchYEMDzbdTe+zJry1+2mx0JcNdsvvkCAA4H2JIC1
9UDX7cqrr8hZ1ty3SyQ8pYjF5TaDpT6LRa6txv/TSjKqsVEotGndnyjYYCqqgJfCb9eZkqQH3cl8
ssf4RWApH4eKd1J6QxiuTNcuzU+5CFkZoqeby+9A088YDSJ3dTRVObRRxnx+BLYpIjtUOOrqC3O7
DktfeGMVuak7AzGH/ICLWsgHgoC2u5DNOgCG0KiaoizlcJlyJU1nfeSd2vjWBanzC0FYq4cCsA/4
YpxK+XOdOAiB4jal3dsveg3Ft2h9xbEkFZBDvcyftJ71D3/EUT4DsohiXubdZkcUqyXE0ffOmT/1
Hw4l+zEN1mg9EWAMQwxTeBQVkkZkC1Z9pR6iK6FmauwScNxGjh/YsNvQzX7eJDb4W9OB0YMT3bFp
zJUK+Y+WpWBSES+MxcCdo7CIFGL0vIelgU0L6au+3QnRmU/gwZGxTqJ2h+RcROtjRvAIxH7iK8Si
gK5r1RLUemRupvlcTOhMMjHJ0XBW/thEsVEkMErnsaYsNdHnBeA9Un1JL6H3dmi3VgRAlJp1YpIy
dDm8C9GPbgKLHce3IS/YcKXOuz4RfYW1p5lrWEQtIBEyI0NICM7WSpgTF0aGMPlvxoWK2ol1IyLW
NnvzGE3+R9HbEwefNC/JCX7qeKZ7wJSZMnUdFCM2Jijetvqu/QDHa2qadcJ9IMEIlaY+MpqpIUzH
RKODxOhZc4wVcZgzgh4o2/szKOJXWI7OZtuCG6WNIAH134Qo+gG+qozRlSOl3rol0vaYkuofOzhZ
YpU1SvWNvp7MN+8DQYfGemmRvGaT2z2OEIdAM2/0SBPk5MZR2HAjYFwVYCR9y96aqwALV8Yx6YAc
yZmLfcvo9yEbOiHmxq8nPB/3eBSZmyHQUmymESl+I+YDE/+Gc2i4QbQpV8+QJJSYAWjna8gDrdXl
XQJGsJ8LRz5xRali4XDeUWMDRY0fGhiLTE4OFbRuAFUc8gVrCecsYdjQ8pcJdOPHqXXRFMXD/nNl
fS4UsdGEaRezJ4J4MrciufXhPrGp5o7nt2DqYW/zwIqBMVJVddyZ0/tC3+nkg+D+ww71j7N89VSm
exO7Dau4HSiGYsMwpWAM88FkXuysPJf/wbRGIoSP1IVZ4zaqLXxUGWXCPOXv2mdfEDtMGniGUnjf
jPcmWYMXL6Y+T/YUD3iKRSHGXrjZDtStJFovG0XYyoh8GQDrr3p+J9AERJU+plL2bFX0vxSGleIz
X7E5+NnrBb7DDljBUwiz9S8s6Zxm0XwmfM+l+w78uFvsd/Elf7eN+1qzpfcqTnaCrxEVc3GY2YLR
dwoCGA0GjdRXISQmKadHJAD85LQ9+AXW3kcXyFgSY3lMturshmCPxgB4scwchDEmcCbDrwuZJ0/n
hGGuVRls5qniN4IfH24RZbEjVcbn7R5Mky1IOebzRjc6sBuK0PzseLWDHPKDtaBdKFJr+TMuiRt8
9Ixpt9m12VbNeUloR65Z1mT1f509MMazfdta94gTPu7xz48+zBKA7/1s5cQU1FtQs8sA0WZ5a41o
vsnX755IstSWWhM2olDvoaTiTvI0SW20TCCHkelxZYBrLRap+2aIPBBruo6PrG1ED76zVb0oaEh6
eaSDAo6iqRhyN60HsLaGazCPgvB2Zmz1v89Rg75i2pdm6xWGg8tzLqGjMSMMVx/ivVBaeNVNpZD9
ocy1cKQKLSChhRYf6yedepC4blG4T+ZryndmdZFoAWu/5ktSrgGaRUAOvF01Ug/foYoQnzq2Mvvr
nBHHQ1GYZHtVCNTJs4XktslsJs6I4ou1z6V0WEhVqLvcVh+J/G43lWLhJV3je2Gh/zUkYTi2Tzlq
GQ0mnyUQ+TjxpTPM4IV9QmT/KKn/Eo+1DYqFklTK9rJK/s7EJBjtvJN044plsZ6T5L4+bnGqfE2d
qCE3Hart2JObaiW33KuWUGVtvsBE7+8yM5L13/eT5TSHmoupaoBYW1FCQ+AGTi66UZZsd82jvdqA
QXGQW4YYM1+XFGLTGuquo9RoSer2jFWorOodVS7HMtgVQFzAA0zK7wY/326nlI/Z+UxBbiFQ65T3
UNJ680Ros7aLUFXvZMLa22Kh2CoJkC+2ivobuw1np3BpYxF8omN1QD/Et+6vi4t7nuoa1L+xAYTX
AcF4BqHs1606hscgmkAHJrYF/4tKxa8+X1PGcI2OfO7slVse51hfq4HhTjlVETDr2cZrqY1JctAt
GYhgRJDbwE54ftKpO7Zbm9T71hSlQPPdNHKTWc/J6HXgP45lryCwRielHmyR2Wt+RXcFXg0wSde4
gm6mCQJo7VMY8t514qiF2PRs0y+1U5AoPFH5eg9SOX+HgqLKQ1LN5LEOnRwbSVULxkqf+mXrSOuG
I+PgF6KekDBoSHk4LDc9Hhjqkz44iU1zbF2vjzWpeTadADsh4VLlHa/jsWpuB6MG1iuCnoUKq4jV
goYyr5kSsq1jJsEfzlqiclwwYzPNsfy7ahRNFcljIp7NaJQ4oyoiTgSk2faL8p6ALl28WxJpQNdY
SRuK2mCtDPdcz+cv5I56rdlyDZSaH35ZjB8uMxgLtf7YBAhv/WAVorY7cZTAWcTfWEuJEyA8Io/F
3LAFkPDcds86+688f4L1P0XRG3YUuAPTB+edDh5yGUexASq3fKZlEXgM1dVwZUpqER5DgiAcMCWn
56vOj2bDGxws5xl56U1ZY5cZSHba1QarIKgwDjSeT0fTLQjYbrwixieuADEk+KYWyg5sATSwrNZA
CQNcKHEGfq712CyqhvLFkmtWUMLN0Fi30IDaFJ1uQr35ldDM1LcW57MTZ3HMg8mC050VipmTL73A
k2mDm9Ej7j/MALpSZX4oEuFUUirvSYAcFQfV72uoyi9IJobJ1F807uSk4FM9hzYjlYXf03ZTsVko
vYv1O/1F5PZXl2WPFt/V/0hk1Z5wv1wHZipLX8qRmByZCA4+qyyfy0ZEUcEzqyeTg2JV1jcJA2nk
5N4jUCx/rOjxwhoHxU7Qum6B+u//gBEL825pCrM0eLrHTC1KRO7+s/NgotGm//zFf7xyXxPI240P
SBr61EWuJmxi3fbmzrgHm/lgzPP0E6zt9hFVDg4JcsUujAO110AqkKQOcfbFWlYlMfS6pzXeR6Y3
/0AJebNQaam+L0v5avC91N83DMfWXeeYRiS3NaywANtBpK31f4x6lVWLVHdUkhiVa5V6J8SvTbOc
K58UNcnEOXHPfdcKWbg/hXNrBPHgbBr0dy6g6ij8ZdiRHfUGnD+kQbvGl7TUE5QqnbsnYJvpZZQF
p6CMu12AIc26+3JSv7QMixtPJP+2KXsZPKZLUVllM+ZyTaOyxBDV5g6qEJFCDJXM8quvVsOOKDhP
1GHkoW6L/GEQwHct5p2T1zlg6ojACJNfe01SatoTCTfHoGdAjDPxORREFzZ0es04OoEfbYAEHpA4
UnVxURyrDudDGX12Wiv/+hXRRD/h5KysiqbRIbIG1tH42S7JBAwfs4Cv5xGNV3juiXPWOaOxi1US
cKaWMZFMDdn68r2B9OVEcXdk51O8+RWsDuMPy+KgG5t9FNpyaABDSFS0BpY60UoDFISjGTz4iKwC
t6JR5TOvZ6zc3yOtFkg58Anwu4sCYHz7qNvqjIGjajyfZ8F8Z2msIPhFQEhauGPWJkemJI8LJurC
RrULEGkLUnixAO2T7j11Zaz0z3rKWypKV53gRGIBI3yFjbQ0ivKbYiUQ1nZtb6GxRvqsP+QiC1OB
zH4mlBuxiRwYkUaLjpa2X11YxgL662XElxV78FFSOilrfuR2L4xWm3RpUEQKWFQ+6yx+VzHcHtB2
pwvdKNgAY4MA1dYjzPQb+GqHl1hpvuxgb3emB1of3HWb3lgnQcDn+cZ4izjHgD1KKYPlVZYR/VUN
hXsh7YD1XFA0CbJtd8CZeQcxtBH5y7jDM7C4FXerNz5iQ5BIOCLBd/gr0Zibif3OGf74/s3K5B8v
1IubssUBHmgUCFofS7jHqVPcnU5RBczScmJFr1N66KmqeiKdl+mRRzE8iTJ8ic2pwX//mdpgz0jD
wOmdiNoyfGtO7RMwVMu0XEilaK0u8hFEPKX7jP1aeIdxOcXfGlOrt1JMMsre+/yGexKVwy7Y7b5c
gqd+mANhbax2RTCuiZ1dshxBQSXgupLPsxtYF5hX2iUGnahCkFqrYY9M6x5Z1WIdO7jVovBsuAcI
diPg3jfDmjthB2+B8gOtg/dsmDOHF5dNOp+TRoC716e+YrFv39/TkQBNq41VjVTqVE9nPpaCFVrA
VQuUPCojiGBaR6Gvi0X44VKp2+zWvsS9jH6ByeuKGrKnhiKN7ydX3qzC2nAYeLO5k2xrCY6ueaDV
q2XaljAjE0DZCczv6n90KJxbntqfSDoqQzdlfDhUdDZG7VYn0zI4NoMQ6rnMbfHv01akrbKMrV0p
mtOlvxX5goVE3gEWPSomN0/XV6KSnu+gzlksXbVvv0mCIb2HNnpVvuDwT1DG2NAvnjww6mZbwoX7
sKoWr01xcWOZpT1/HGRmBQZI2EL2+s2AZ8+QPoC0i2aQPBUnrIp/4ikUE0KUrheVX1qvPlEE525V
StRyYTUhXng55dgY6//kggoJoDqTYJWWehbEd2OsEwwDb5e3GdQrh8xo/kBrTLdMxnDGpG8xlxe2
grIyrjvB59cpm3Ct0TDLcHr4pT6zH64AbtxnuF8lPAeSAlCnbQpS8IWbnU7p46khNjkSIrQalivr
jY2Jjl6BSGWrw+6QXcAP+9Fb5+4d9oREOTrbU2yCuFZJexl7zA1XBD41DEKZ2vXIkvdhhHA1arRL
qKC3czNTN/qfoUPybzARFDv3S8wfb46ZyaqDtjIoq4okpUS1LhDiK3l4Blr+WJKUJxlwjvq2Uc9d
wKGUroBEMUyqG3Y2+mTB7++Oh2/imfjmkRmQHoMPHoE4BBiJ6l/8udEMgJ6mt0dbQjlheeSCr95K
1Z8LyPtmCzQGMNqTiTEH6cmGwhx/zB9y20siO5cdJ3epo1Q2KH4p9kVka4TIxafV1S5l6+btpkkI
QkP7bErr4/j2Uf7LveTnbtZOdeWZFP7tGmkL7q5ftX8fsWg6wVBZlOymei43w4eWt9WtTY9BcT6I
t5QwgA4KaSLlSFxpJkLBPMl7IHa2+Mo4uYiTwfB/aWMXFrC9s9t2A/13e2WNyFworSCw1GUOdQbR
7VSAC95KZgfVY++YofusnJfkCYyjf6qN30soHgwQJm4aswfC89HadFfduwrC6hnqf0N2t+KfS35p
VRlqIX+ra4YDKO74JTSCJzi76f082CzEjxfOHDtiUpTSHc7CIlonRFGOw9hRETIPCsr+R4ct7Rij
fgwl5UMfge+dEI3Y/hSSTL5IHWFBfN1dogbUTf6gBbU/DblA15fS1R5mMJ3QVStrZ+ZbeX/7DVJC
TVY4+TkUpBBlKM80IEGs/O4q0SxpR+vzFcQoEtXBJ55577lXG1Pb/5GrBOxBgK9gvqelFduw+mR6
SyJGrq/qirENWz5yJ/AJG1DeD3maIFuTzLqdzdB+rD9SGxC6xKSiFp6elPlc+FqUsf5Pg2XLoBZT
V6Q5G+14Ex0oVhI29datvFR78uaiB7lhJPp6Nz9/o87HlT/yr6rhYaGYyzWdDtMY/tFaGbJa/ksF
fW7wROMrWyZ8F6xPHruPLhVKDD0oWeMeaOnHfIAOeD1+JJ6LtA83gkmZ4m62mbdW+xVEQGkoom6h
yHqna+DdrrVa9RpgeBAhRmgY/JtefKwl0viRo0ZnaVl1TpL+s6nAnQW69yBMO/0xPm0vPA2TN+PB
01wCfsSpAYUmHOp5vA+biGZcDPOziv3ER0vaz3j/tkmg0ffstHlOkZq6PH8nvVz+SGllAfVk9axc
//n9zcs47MevuvIb/BB/PPDN39i88CrtQ7dBYlujrwmAF3HQJ8Pac+FrDOGMIpojThrySw7Q7poU
ve7J71jUF1+7c5UzO48Qs/c+z9k0vUAvF3lF6nZXKpUIyOYY73t1uGYEuqsTvsvorpBI6XyIkpmw
EScMOOt0HXFFJlrWRNaess94hSKCDrmb1kN07hRfe4PorIxWManjCPEf1Kef/8IWqPdOiUILtGow
E787WZBJo9YsLfkggMaAXvvvVNceKjMUDt4qwygReoZZLv5OPw0WP+voZSOIzJ1dMmAnqgJqVVd0
/38/30JfHf19DVCZdBHbQguFpTQSfVmlVollR28vemYEEwsE2rEH2AU43HF8JMsoq5vzod1cgUML
bN37WSIfb6UZnKXTe3392gRNfY5VTO4dZ0uG1TN0apVDZxbMUbnWU2T5YhLVkWMAVV28RN2smwZk
Aj5cqVsQh8hYLGDZ81xpj1i39PePSFflVIIvEJUlRu/lSkM2NAyBZ3ANTkYUVkUwab6AvvGhfNwq
SS3MVVLg9x5ZD/BqZpvyQ7ANxl6fWur0MlLGRHPgrIlBkzPhH5IGSLSkem2ujHdrxHPjV91bMOh5
0e4FhFobugukOy7sd0hlDgc4jo0jUrwhHIJq/4h7HC0oNeidrccOmORrxYvBrpDhxQcEgXpvsDjq
cwtNkdZhmVvcw6rVHoV7y7VXY56wTLVgMVq5THwB6oQjJb1CoyJ+B4RpCe1cb9FXoK1a/N4K9vBZ
AuvF/nYWXo8zoBjus8qtLvuWXwxzA2jQD9HIXo91vJwgzYAjNsX0VlKEJcmubtfgKk7YZl8kgaYb
n1DNuFJTOfFCVOeEOIzShAlXi5rGOWtCV67lr0s5tf4z+WU67t0JXVm2eXpZX8y76xdFVOcJ4Uvy
HsAjGWGNW0ifbt6lBT7R/btw6mqFSLFUhqMWRWB00Zy2mQrBdvjwMyPkF+ps6wVd9N2viNUVDDhw
FVoFou2Vq4qJ47xOhvXhPK28imccRMnR46CF8jYprrZRc0EFvJneYdbG3OdwZDICJt7fZtWPi8tn
1plwT19Em+VpgSxFvpy+VcXkualhA5evz3nVTbUi96HhS8L0TWjrnqeHEkYSq5xKbCguV8wR1cBQ
/TlZSDKDzTASrRXgn8m/dqMNq0vIykghLqn1uZEK4b6LXE3bn0wox/SXEw0YY+w0Cwm+N9mJONwu
XXtkDTr/pdY0jmsT3HcXPY5SajZ7rz63NaV2G8Q4x45xl92IGtbT/syRp+TzXt9Yju3c5Cx5OeaP
A23+haFufVkuz5ykuG2XFDlDFZwB2b5G3eQFa2/46t9Fdnpwb/nxDNpmYbTrmcn6Y6n/H+iiqO1Y
iA8z1x2bVidzq1mqvkatPWHap1vRrf9e8w1UCV8aMHf1DurV9i+N0r03hwsONEZ63QKXLpUlvU4W
49/bMwC3oaBTM8fKiZMTKYQz9VnD5TF4YH6bGlO8bf0pHThCxAKVZKWH6Yt04UDfrb/hnYsV4Vcs
2JKXTmXKRgWR9ss3j90OjmHxm3H49oQ9hqkawtqY+mUSAyEW46B8o/6WIA/0nqz3V//UzOz02VKD
pG/4LS7HQ2JIVwI6oF8R55+FOkxpoglk7jj7iWUwejZlMH04KKBxowxtj9F9tRcna7+zQn4aqmVq
grjNmlIdo2IqgrR+UWg9ydP0XY73jVgghyaxktoDU22+9YIZwCbpB/u4FN4xqBiwM9l0TdO8czBE
yV1+pFdTiyvNWEl3Oxx+b98p+NHBmQgarU0k6gm+Y5+5/Ef9Y5CjOrOOxyGLHOOJbf6CTJvC0wPO
GxITWX3C8cT7479FprhJAPnfHTyWmhzW+25SpW6KiF9cP71Dp6KRxqDbAQTMVHNehnLKTf5RVQRe
YID84O4TUJknDuLu3fC8uz9sSzqiKoVyppB+Yq67ddPU2kE57WGLoAUGWR/6BDAwfte4B27Lr336
8b72V/WXs8PiqvtPubcB7JvXfvwSWluABwOghGyHgZ9OpwUlspuE4PWdpLS+XbOyWo6pgKDoqi34
dXMajpEajlK6TKLJjfkxsX0wrqQ4HmNxe2pQC4Zih0VDxmSw9jC6CsPb5bfJWmFoylGRBW4jjv9D
XMJBMfpaO/A/zbX7r4n/+DK211qPtmHovK5BtEOfPSE/YIZ9pK9uHLdPsfLRXqJeXp//9zrm5kkt
ekr2G7qG7io9Pt+BSqQp0cFCffD4PCm7zC3OeXFO32izursroplbJp2lGu2ARhu6bvTCoiE5s/L0
HoUzBlx5boz3XqlHj2vOFJn0h0lIIC9usw2OCnWNpgzwBNeo5JBt/w7TMZ9ShAbGsp2lziy3Hana
63UyrEKCYfNHTlipBUsOGZO4VixJyMwHd7xlAgtvK9irgaJpl87TdT4OrlATxpv01Rb0W/gp0hsF
rOgYO14G3lVcHg6reHFtMaTYNQ0rDCXh3ihZsHAam/KjCrreSmYNeI3Jzmwkmx+mx1FZY4XJ5+wQ
jl/kz7ucs1Gg0zbLtl2NjEyvEvgK2+VXJTs4R94PDB5zw4xPWWFxG1rRGu2Eet+6DVd/8qLuVKax
XXEIaDpOjVmhOAVLpAYOG5a8Yv2QZnZaAk3Fa6inEW2INSzuZ6Svs+lcrCnN6rf5ChfXZnF+aMQg
klu116TxOwGxk3H4nlCuThABzVpSlNk31Rihdr4GOGNMVeDWj4RP+xXiALGyJiFxF/E2dxtFFh0G
eoUPPapP3NSw8m19yIrkMQl8lpr6+2f2rDVuBgSQ2tWZ4EEtrcdhtA2E0UIMmczLznE82ddX3bIb
6xS0ces7bU0h24ZB7QmXZ+M4jxNOxGYSG350nT2afnZQClairA/TNeGDpUz60zKVuyNFeCPKUBrE
+5aPxwDUzwg9y+i/v+E5iPxURKzyLdWvbINSCOa/6qA+m+mMjMshWDx37eaA9mhPf0CMOcpantHi
DgP7bnWZPhMcX0HCE5gOu9sk/7nHj574keEJk8KfnHhkFFyuxUtVppIZCpyojvmaNMZUICkM98rf
2fyJOaKPu9J06FnJLD1Vu0mdxIBOpGD35OGxdLD3M+tRdF9ouBer/cywydDeiMdz/+mLutq0h48z
bWpDzBnsIMW/aCoeFVpwJEwpWIdNbl1CcfhtOlxKfJaqlSRNYK9J08xzrnCKdpu9wAVl5YoCyGxO
x3QAna+wvjZzk7eVNhXu4tXjFy/3+xJ3ee6MyrG8Blym0M0PRm9Feo/jPVE0KRfK265pCDArDmKV
pipzuzDLYknNa9+xnqhWUOEEKAJmqZtE8m3/xgRGf6f9oifTX8EMQVXgdX66MHS42cZzJ/szejeW
uq7UKTX6QDOUHFfj7dDelTSJtXUGjtPeczL+QEopq1v8gPfwe3plQPPOmbPeIkvfxvzQEZYVCAXt
lWxgl0JMhNMPSK7TxBhi/AwQdkFYhtkju7VBGUnAU23E48iNqIDDHfZ4jRIafa4vcyjt6JKBdwqN
ulpX+M/2Ws86Y2WsoziDg2yOpcB6xw2jfwMDwva0uH+GxqpuwmZw/fhY2NSvvQRFTCtwiN9xRmHi
h4ngmfNh2TGrvN/4PPFCuW8mMsrU+qEMmO6GG8dUG/YwBQAuCiLyNRyOIF+xAq6v2m//8Tuc97rd
neSA6RGLkllYc61I5WKBskwcUVF0cvBTALxZeNjUMBV/FuHaLoOvlbv2Ey2QuR/65Tr574lFPZ6t
InIAX6cvzSDp6yLuynAkpAgzgIjIVB7lw+mfmQNBqJ+ZzsVIqCb2MXMMwwnXZH0h3E0kkF5tPNwc
yA3tAvEVcWhaK6d4DF8EY1qLwQEZLMZ6Qbl2BhjIDrdwzQ/DM25VNbLETv9RnW7s/qNdxcD5TjLS
7KCK8NMXDR3t/RRWd3bf8xa5mVSFJSr9nitu3udVhVuv3kqlrRAWeKf2g7GPdJTfRMYXVgzBbTmn
+j9dq96C+Ho+ktKK8Kz8XUlle23MvlxjAr9h/0QYa0uo751cVRdAtiz0TkN27gdaCJ+ND8552MMx
MXd/x1dzIddxpeeYJKSPN3D6aqDYYoq7Sixy3uPccTtEAREL/u9tVc2nNpvUUxsFrb5X5HZvWn5X
WHvuaIHYHzqRybq5OZAjOus7JDLa4DwZBDTNQCeonB7u602arORWWeZ2AcOrPXV62G6SQgJfOHml
DVGhcexeozwM0HAUGrFUBSXth5Y62zMRrDXt4p9+JufaGrjbbkljkdEj3yAfjHak108pT/U/TDeI
G7idsl/VyGm/b6HoXIRfesayUUbt7+RZtbRXusoXYEgUhCiSeHdFkOqnrvlDizVTplrezWyXFYGH
znwUChSoW66xHipPVQBh7weGkGaX6D6bBDsA2Lhya9fu6p9d/R/VQQnr7ZGRWQWJzb031XnS5raa
TQfSLDycyNS+ZAe3x0ydb5pOCYdaU45tcIL2uQSjaWMFxUzrxRkrdmBMGw40A5lHNfQgcSIxcrM5
VCXAkALeikvA156/OoW1YmfFF0mqyVW7QIs5tBl6GUJVXnMSQdzo8qelqPuwZn0f/vTixEowW5RI
K9+GwO1X2HTe8tmnPy0m3OJ9wfnHm6kDcssxNbTaig+7J4/wVX1PP/m3iSCExMCmVekDZYr9WAUJ
9K3R9dToqjHb8R/n2KuopreE+cwiRi2XB6clk3eOFuPaAG6qWzTBXR4VbSrLPlOiIvhyWZcw3NEf
qp6C4kCsWznfRMBwoixgIt9oP5aU1V3WTrJ4Bvd5rsxJ3jDEPtqbHRuaTxA82pbuAyh74NT7a9rx
uybZX+Y92Z6DGuBGK82iNR3jKes7ZvNIil1aADNhS4rY/O9Q2WDtFrzqs033hLhcTvafpcaEI9a4
7kHq2QSPqzzpW6XAcW/9eRw2K7gnDi8QJihy0Z40USz2CjBZlxJ7fj22JkwUp+/tvphPIKvftJnV
H8VcAzhIB8xFaiFqmk1FezWJtgYQ8r1aMYrwsMlz3tPJjXtV5fwrie0NpGrtQ8YuGRDMi6m014JY
LJ4LsjM0MmKwdft9q2aY39FJwMfd/v/dAf3IFRzxAW7MjTNLMsfyk3kx5CmCF2FHcszFKKWy9E9p
N72jE0c+hv7cQ2J3lMkUFlVhjRcYU1AZ0LstGxGKZvnJUnU1B1tcsi274dOWD843ln/FU1H+Dehk
NG7zGizkIjxqpMYXAm6ASyPhkat5kgpHOkcbWn6KtBaKJh0ypOPhqHgHHjX5cfjR8PElHdgr93lQ
4HE+x3LfMU6sM+Cg96jRxcgD7OBoopzSBh9b5edlqSekyHTEdhbQlyWqjgZdwYwFmSIPkVcIKrGp
iyjHgCvAki2zw2kjyZxAICL23uh+jW6SK4fpoEvitUBlB8Ez44jZYNXOoDdqf+PIaEy3zWKAZxnl
QA+xTNYCY8r8444hDm9AG8T+FWxy7I8rMeV4R11LrtoBZ0k/wonMElETEBYbA9JMlXwxgPFWIfRf
xVzb2bg5p5HWBFr1bPMouzcw4gEN8bzDVhk+qJN+aiZU3v8FQSRt+pcjQ9Dr1wULYOJ5vCWMSBK4
sGMkUWM/AmgbOZ/i/MOcl8Fppwp5djZ6Ub2Pheag2MNedAVlFTZWcPpGbUzSIfcLCJRGZSHdengD
VReJtxBW/bVL4P0dpsrQKQ3+cs0QkVvpLivTz/lQmTv3/AVNJTWFqOneWNd1qwgd5WiwEvNUXUO7
coqaqvMik1kIUL0IVEeZwiF5bbRUz/XNaZ3dQHImjxlfZZ1oJqXM2O5hb881YnlCF/lDXJzboBDT
IlPrsGajEs/n/cXsGMXlIgzvvQhjcgEUMrNFDImq2VIjNHEFT3QkmxN0OP4xHWcQ1P7l6uX1RC2m
FGHXGSYYafN69OziZBCqWUSxe56BeHU6aDqGxP/GUndWLewuBt+yCRfGagWjTEZEuz235u32UPEy
yTXt/e27xfPj9LCFwb7pq8aGwMRtmjp3hbFZfFPpazBsFj/LL/azlu/r64s4Sq/15eIbml5COlNW
ULwqRoOYCq5s92/DKwpJLfXHDX01bfp2owNuySej1e76pFUdVE4ITj53ZRJ2VMZkA1OyOm55WLX5
xD4+d5EsGsR4DKs0jqQjdrWWlep/fDCtzv1gAiAky/cqJoZIGyKx/IrJHxReYAGZG4lrAO+jU4xL
s4nXhBfSAiWLdn309TqBkeZ2EDF2C5F835QH6udnWxW+7sYOFv5SpdoYfDqvQ86BjeYntjfcJoQv
m64CJThV0Sr5xm6nh2E3ZeYrgSjIJhLIeB20VRKtyrI4TYARG8epZLjCkoDpa4j5RcPK8l4mLJC7
pAIlxtHEJunPv4VrSIt9CTr/8eDPcaHY7cvEZPUPw8Cr6fIkQ0/lcHYLrtiIpck0zQ50x+Q4rNrh
Of8tWwFQz8303Z9P6vTx1E5H9TH0qjs4//bgJIt1clcmd+6uK1l98mabNtsSqRysS5gaWY/OfoZ/
RGVwU7CU7agJhjXq6Qk1pUVAqr5AJ8bVafbu5qOEAtOBgW/iQWMZFwDo2+Ofes0naDbGSJECf77o
/O8KDT2iLd8b1rmfuNn+2bG4Y0iHg+5XikBQM917pIEstBgzJRwQnvdmCNxN4FbU0dKXL+v1KPxB
k41Ff+UdKbbUyS9og43WlrzWQ0elU6tq+sQixuKwCHXqJIP6HMCa9QQ38WX8HUkQrN3gRKCKZHai
l00v3INfeZWp5Ev5Ku5n6+MMSsIMrDyWvVTR0pflYryAEVFiPluKGFFUQk2e9cdjc9Bf4QzWHaZp
mjA5UOKlEoOg5sbO86fJaRbNqaaHTjTG/8v3FDaTcFaUFWoyMjsRlXSP2aSXJC//7vTwtssC0Fxg
NZdlbrG9mxDZ9y+MG76gQc/tChH2VsaLfGuwM0IsPaz9R16mzzh75H7gjtp6RD8S8W2nmnOMAJWE
K29cZBYmcxONtLdqEWT/AA/Vx06EyQ0WB5zNTdwnrBeqoHXiz3x3YLBgNMDXSlgfL3bzVPOlkieO
ED4Pn76uUdQ2QqP1cJjZxWAL6SjWP7ZeCSj4sU7NtTbJxyqU/WxwdMk7Mv+6peq0nTyVYXZcwCnG
6ChqIH6T0gs+Pq5H0jai8GDw3iVoag92nihWamuzCwGO6K/DN3kuhzl7HAe/dbUiP1vsd1pNVdMU
J2etfA+tf+KcPz8YJbsgqbvDrJr7kjmBuw1i1LY6bzcpwiWqZIEkJhnO3l3jXnZEWypHxrNQRYqE
X3djegBNHQX3JVB/djIdu7M8U/mLNdJQxbQKDmItkJCD6LOiuIx987tC55M3TtERpLvBGPgX4Tq0
s1w+XZR6osWqCj/1PDbueGk1yfCIifhiupE/0i/t7bCGePa64Tmx1KKxb/O3VxxSGM43sgmzxEKY
LZ6UsFrCrVmKqYTgauT5bn46uziIWgfm320Qzr1B7v3P6GAFe/T7VHaF4y4WAe9mcCoN7MENefmx
WT2gzXtHi2U5TJo55asetJSGPvubG8zJh/03MftbpgNqYoT+82hJhmz1sc7nc+TXqaDj1QRdGVWu
yIt1TmCvOwwn0AsW1NDWwS1ugjUa9tm2ryOokn2SI8Wu3mdi1vFOkQzdwItBFvTStaBoo85mcoto
jHUA4F890FiP9qzj/8NpNj8FOzxd3+ZSzxvlmfkKJ+tfqcIjZOAkvq+hODgO2IknViW0Mb+RRZ+J
/WjFgIVwqBVgBkVFPtXaj5u8028ZKAJnUQLJXoJhloOw0O8nPtipKmS/l4sxWHKW2kpRroFkxIJ8
wYzm5kQEjRsLmP9makTUWk8Ptc+hS4ExjA1bOaSJ/RfVRoDr4fO5rQKcxyHqqHTogS4gzjRQHQ17
xSg8AsEX3N5GtZjVTBs5yi2bkLsPIF0uuBR54Lmh8C0mxk8jfeeN65eVMwO5KlG9iZNhP9D27gjg
bHTPJvaLGMZj02G9G7m0HZk6atVnnDy6Du/FkeKkrnRVu4ufh5xIL99q/k4DOnARfvoXd7kpPNh3
3sqHFxF5CY8Q7ZK5eaf/ULJoBqqbAlVLvp+C3r/4HY/8eccVdlHrxYtvhUtjQ6J3rw6fgrwhHp3S
Ex802GWyRQentLc4G3I35WFoHGGHkPli7oPAQ8g8WI/hZ8FnZ81OAfVKbk7i8IFMa043QeoNA60q
yo9+QMHIhCWd70u3nvIRgv5oektWfUz36DIwIvTqCii8jxzBBeN6EKXceiH8Z7b33aMAoUOdcc+I
tTFoTDbdEvVNjix0EHF+RXKAjeQHEIvjoBJK6MtcWJifgwxL5C1QY3SlRuZGZeg5kwfPMdw4eT/7
WLxBdXrgvgJfRNA2Y7S5CFLUcMaE7nr2AmKai9jSetZ9GhNmqYI0YgupBvNDfH5R6yhDM2/alWvg
aMZXvTJNJ1WIN/YuNys5EEyKKJA6UY4EIS0px8sZU6zkjM3tifLrXlhKjJ+IKgBUU4lzClrqOOPx
fJP3ftLyYUMshWFX/84UEgrNfQH1ESPbxRYFg4EcpVCByptTcC+vAUKeMqbHSSrpvE3ug58Ubapt
lwix3eRmfeSAttPqxkno5WCNhnA4OAlbXUpplvVtYDIrwvXUWbqaJos4S0eQfr3B1ZULMDbbWSav
h+NnhEUsRLZlBefc75sab4COEik9iqHC3l36O76bV2A1DfEA/NUF4ikdp8ELQsu1TCECJb2hEQwp
yh3unyZ6+3OF94zPsL3JL1xK7aIvgPOoqbuwf4cb++YBgNpcs7XEtQgTmlbrLh/CqOumVFTQasKD
rP8/Nxh8tYzCZBowWYZih6G0rAQbncM4bvD2g2aJCVFIlY26bJ5oeVNdD/WB3jaQM0Qalu8/PF9w
qsjQAkurH/DLZ50MRDkRjSz45iDoSmKZVKPme5yllLdYMKPQesQ5JCli1kssIlo9jWjgwo2xfqQj
ccVxjUMBWlXa/sKIvtdhOARxNrWGKZTRPPruFIyKG9gZzKRVPIVUE97LLkFuvasbbPglhecinct/
rQ6lF3DMZ/GvUef409ifIn89ooSkQOha/HQ59UyYdl57IkMGokdKa70MzQ2Qk5pXuYtugrNjK0Ys
KJ1K2dXxax7lo/EoXP97jRKZVDJqCP6koQy8bqn5Aj/daPeVLJ5W16v8UIhnG7riNR0QSMqtTP0/
BMe4wOcQ/qlRRXpUX1oErfNN2HPrZzEoyHrJi/6xX49Hr3unj8vwlij1WD+dOknwib6Shj9+HGpe
OgCwDZZ2dBJSdlVECHNXrKnN82L2QOzfntETBwKKg2RddLJ7I03Dg2+WIS3JIxKbV5y/HPdT/LQ3
9HuKaWfDR+2nbwMyPVx0WreRLiFPEoi028y5bSA7ttuloIhV+bkO0X2JVIf9h3Naad/yCV7OahFX
24dCNEm6z+uQGJ1Dv4MO9aJBNgOLtnqy9M0LC9WcQQ0C9eI9Ky2ueIk/QL1bQlDSblekPVjUwFW8
mzFjXU7cGweRaxwqD2l0fJyPl8fItUsPTKu5f9qLC5Reis6EjJZk/iuqWmxMPUHxLmQeNNMT4avZ
lSjTNs1GOZCzQ51rMloMfimlJVLFJ5L55l4MuQSI3mvocm/sZ9QnqiYSHRnloyT5m/PWWrPNuI8Q
+f4j2c3biONrZEEBl9tLwzhfdovXNzyApY1FUcusGgl7Jf65k2a45IkD//z9EqDOWgsxryOX2JFI
gq/oXL47B+CuHKLEjelLVjZgmXm8l2hSV1Ph5h0q5WUjK2+kMbeXq8gL9cxfxYn1B0x3bbqae1KC
P1buuYKzuAIfT+hf16BiCzTd0uQGAVvGDGFy2yecRslPDoxPvwEC9moFkS3/qdY4ZlanRfbs5j1Q
Q4sBKpzS6tpRM93NUluIhzoAJ1auQaibGj1uXJjo/x9vpsPuwo7K7dlDAj0JunRX+I6Pivq33rk4
Izh9wl83hd+/TYQYWiVJkOxM3QKd4WUc2CkPPY3Je0TzRo1rBFxNx/kCz6YY2o9MZwOv7NA7Yxjg
bjK6qPugsTdD37lgm1qeygwp6N+AFU/4uzLFJKC+1lcz0UjnsSdcOAO/LBMa8GIKS8ZZLPABLea7
ejKyyR2dIZ97dnXSbTxQ/ui8l8NB6inNSZX5KcCPHDKn2JCMomazNqU8hnlVdN/SpVuzFRXeig+S
p8LoOZAoNs5TuKzxPHtKBbE8cOPlJCjaKrXG5l09Am2u9dVGNge9c/OGxdxFKQRaFlSy+QCGDdz2
zCsp3W2VCT8R12hxUm5UOoAO184InpspjU3PiC3A5qFJxYAdXgQ1hQf4awyXmAn+ZoOSsMmWruyT
u2xocNRcNuxFGly5WO60fno6e/fkWyI6lTn1dby1hGzmfwu0GZbVkKi4WMMWO2LzwmqapP2hWBbi
FpnURRkbQjJwdFrZmYCqQ/hikY9m95FzxgC5huqSqODi770pJ77m6yiDDHa7o5ssgUJQ0k67iqg5
tmTrOSz1TWYVB3mZxzYHUG6i/nRFwGMyULfVlkQewww6oiend9Au/iLWGRF6N2Kjmzo9BIEry0Fq
vc3GDFdQsv4iWkgbnAxfTAp5NOGVcM+2TbN5Q1viII+PQudwS0BGBwYxrM5+ePEZwgLoxkQJfho8
tstSjUcXqw496tbGsMtYs5GDuOiRUverQqT8b4zsb/5tlSo44IeUvACYIu3V5bfCnPN1NHY/mkuI
GN13SUPNTQMavXpllbNch8R54Ra/T1UR50w8o9t7JFK4qISqeK2Dc5GUaSPEog/eHmvqVOh2hwWB
grT5mJuY8s7OfErBO3R7SguB9uCaKKXqyn0/RJEuFaNlTt/GJu94SYuxKlnk+irIJYSm0P3wUPVR
OnA7lvjsdD2qt5uzrtNQzz4LKwJzFXwe9fvlIraBrjdn935tCOeZRRC8uv5kHWf4uXzBOozqGvN9
N8BLE4FIiGe3S6Peol3a8Udl/TUo2Z7tZlOdQKrYnVtCcI9tZhoUGH2LnYsX8S4QbQWpK+vbG3m1
wtktvux6LST7/Og6cDidXHEDHouu46juUjK2o8JlJ97Q7l05iHgDXp2LBAuxbkHWB36+eVM1gTXo
NkvONBdvUsRETXgxJNcpzwBXYMqRBEf5BTQQgldQ+Sy/n738AdeDQBsVCOhj6VDclvry2De60ayG
Px02swjSMysi5vi+mtGTH/x5fUX70T6CVXm0392/uy/kwsqP0FtmXQb0olhQZs9Ac3Phn2WtDay3
2blCi5mpwrYg/Ewo7FenSFH8t2JIUlBhQFniyZ1DAQefqtM921U+QYWwvIPpvSakS/83AKdMVJw6
t3WPTLsow6VDKSBbAGhVzSw62l5QfKSgb+IorEXV6XLSlsoAh4ny04FYNSIpPSUZ2QJjbQyAtAFV
YOftxh9T/QQdfGcMWckVdir5NpkuD3k58t9d+3yHR45xA2jGDVrK++pvvEDdeccLKLI/t16Ef5Lk
ZfEsYwT6ye0GnGgSxpyunpY7hRh7Hp7zpveUkTAs9sRqncKpjFnzAJxWbwfy3FkNSv7RU+upszM+
kZHp9mtev7x1n7MTpO90SUoWCv9j2QSpsGgnfkCl4eqtVelx3dYAyFp3r8H+u2vBpUAdLpQFozBB
ozfOMBRuMRm6MWyqv6ghqJIdFidFPcQNZxB7pop0oljbzpYuWtNCu37dxCunXVvjGphD11Qg4VvR
reAEBcvPqRhBT2eX5PKAbYZIQKAog3+Rwf8xEuCJCbjyrHY6a5zmRD3kxKoLCXWKZaJWF+vBJ60h
cZYD/CfZLKCBed67V0ha+yJHqzZZT5v3jhiTAQe34H/dcJvk4t9zhqedCloYL4kexUFV1jq8v39m
W2vpdeMFQsoo0AzLSHw9pdzKaL6CeILnCMEUryhaj8Kda+sNPWQDaF2YyBEUJFoSJqTyG9hnqhEm
ldKrDo7ilnqf2cev3ZrRlBInM6a11FDPT2UQKf3XmWH1nTzlpE6QuicKCWvFwl6q1in6NKPNSYSY
oSS33ss39/xNYc1gpw8OEDt4NKDQQcuBHm7LFQEoJycuHVTmBgCj6HEl5GvC/5hThJ3KEKMDZRff
jHWiYIDGT3QdruE+9DjQK1h+C+Za/NoM8xuFIsUqskBeMfyRnEGU/J3PVg4g7VeC095uVJlIX20+
9RbpL7L40gR0ew/OaBcl3Z69hjZ9rJMZpd2hqPU64ggeGUvqqN9G5J7/yxwinooUC1JzBIEdEVWo
JeQc492IKudgYLS6qHgnehjUo93sWZq1EKM7BuTiAGve8CPIIDt7N98isQrsd3reyKwPxr3Oz1JZ
eJGAHjuFs+VCAgl6SK1Vol47HAiGZ8SoOJHyaxmT4qr832c/+4lslndG/+/BSSIvJvAYRh9IdQj/
VLQgXoBB22XkHFN0YMPAcLndN7tPu9swbFSkHdTqFbywSGMLh9gBXiPIKlABKmjFqVJM6Ubn4DP5
BTrwa/tYXbO3KYex+mlKTND3VaoBMHrHYe0jN07/S00AxmquQhZdQtl12J7shXr1Z9HEVaHuO2Pc
QG16IpM/8ZsjJMRju7U+zhOe/iSyLEcyHZqnwMP/dfhJ5SvTomf+tm6JVDEd7yXHBmVCCGZSenjV
4ph3hHRqzEsROLpLKTQ4l0BEY8j9rURnVm3ycIr+63iNcjHrOPBESdIi1rNaH2EsfZ8bdHiq52Jz
GUABryqTrSAcvuB//266fXWuDvAui9h++R3dHlMDxkhU5BLaJRwtUB72jaWEV5BEC5gHWwkqkgjl
nHIMvMbYn6ryVU5fqOdcyf9z/UNXIWM1XqdnVEFXrK0AfE3jxeW0hxZxndGS6t9YKdRlaBpCQ2pW
7XBXnf6q2SC4Go1JU/0heyoN8OIKoMSwZfLXpuHXIQqHIIwBoqUMVpkzEAC8sT/a1oOiP07GCS0r
u4kgwGgile04ojcp7lgr5NOJy1BBpKhBGfsw55gApKOPwD7HCm368Tz78FLiyLBIeLEQrsSsucNs
mVj2d2Zu8NkCxmUqrzJODOpKnaRq4bZtbMK/nixDaNBx6jcRPbBLIjhouwZwoBr9XTE47Fx34l68
8T1br3wTg9WqMBsKdArjcVSrbkQILNSZIzoPAdvu8owEpIHf46enr8U/poIwy8NSThKKvyRygrur
awsC+54jib9CzhVLcy0PgCsk8O8VRzs6zGkZUAh0V32r5lEXqGn+av5aVXxPOx8I6bgrmKYOdqUZ
ZpDvaa/dTB4rJPw/gRMS1iAJjNQmwV9d8zPiMEaFEGYM1xvNfsvIMdNcRrWa4KfmWh4Tf7Qne14e
VNsL+tqGUBOhpGHTf3XnvLS4wNnytK/4XcOqNxQgri9HMzqzlAYRRDTZPomm4lUK/FGp+UeoZBQ2
PNkCFnm1kZhO9FVB+rWMJ2Zs0QUs+ByCouq8TKwpllqktJN8XwJLQMtplP0iZLboFu4KVvaEg8Mn
sFK9+XqyEr5GX8d8MW9/3D585zcZlpSMDZkJ8doNFXaf1MhE5HgbXW4msG81UyTEARZPK8BAihFV
V99hSrqbnIvj0+P+oaGBFA6KN9fuS5g6qQylgYeYDFGc936+EHpQRYvil29V6htKIRhUgH2vxNVp
SSLFYmci0DpXFvJG4uD5RhsH+jfOwn5Xg/R+wRJWIV457of9huimzkGXCcXmePR2sejIWgSWHV2d
Zn3xH8l57OZbPhOgoXegwuxgT558/dZCEIG9N+cERcrWsLhugwdhrHUWCq63Zdz8EFaIvWAMi/2K
WR0bV3f4A8ResTse5pshmibXGbKuMLQt7p7+wI5o50XYoreg0L0TOa5UiSl0gAita6z7XVTNkInV
sZ3htpfHxitsUkoV9RRphwZvSqeX6HNMEgSY8etkXLxpBIjWCI8YSUnF8oNj0SZ6TQr7YzihU7lm
H+MXEBwhdiqBf4qi6GY5bed2trLQp7p9R+YnuYZ9L/1l7VEkRu6lkYeukFtxy0lo9gcMZvjccMCR
Zthwb4O7GWu0D0POls25J9ZEEhjs6Cs/fcgKC0Jv5r690bgkFvQyJUu8hvd9gzoiZzeo96rxMpDa
ll3wBvMfHayMVrwRL2mcrmufpgda09OmSs/24BpoGioxy4v0R+9ZO+PbWsEifxV3qkVOMqQbMgnz
cDViLNoqhciLvD5p7QNlHCUyv9sO5jypo0ZnBZgUOv6oCgWvgsFG6yicp9EAn45nbMp7kxUPFrnx
Y63/c1FdyWrmeu5xa5HWZTIKll5F3y6vxN1Zzpi08VqbUqanqGa9JHBfVnyi9AOyCep8tjecSCGi
Lv/dnO0b0pry96zX0v1aNOpJypEHcIgjbTzaBT9Ha8EaCGH9aL70pRlWGjVyTn7MIxMcSOPzhd+m
KmlCcHySQc62VDa7Ho6osegIDNoRkPWxhDTl8koLgR82JiGzAynq6Ea4D4oa46Z9x5DGFOC4eOel
VRjYGB08MOYGeFWMVF+VkbBZV9WWjsWRZByQ8MZACizdHwdAk31OPKPQFkEYnotgvcFxb2rFNrwH
AsAtdBhpNDmXvAMzwFBmiyJ0LtAuEceEGtki1px7t8voY9+cOwPvAXdmYio64+CsCL/Lxt5R4hNj
qTt7qrl68NQwinq2wQW3UjfBRbIt/acZTBOhRr5VAvgcMz0p5Pv+1kl6fYFy5+MV3uNgm3Y4Da0q
9Kg2Kd1nFfp6erC1XKLahF21Ngc+6y/JZ+N326M9bv/QPKDKPflVEvRzM10vr1f/2w3iMjdTyA0r
5N/VLCTbVfYGhk8DAMeghKzB2gafzarWiBAow1HYyKlSdGRZbiWJqE3mzpfGrhMhRpxaCDsikqUC
5hpx3b5ooND2y4iHJ0m0uD4ZywPAq04Q6enL2P2YSjEqdwv0ZYmqMDTZRTsEq7hkvKD3Q98uWTb7
xvJbcGOXWqA/jQ5ZwXRxoU2TSqSb7V/fQtnWuYsQE0aWpnyPM8P66Dqii2m686dVlA6vRwUP6GU9
pFdZS/bzQnaO1PcU8soP9mYUlF4Q8RwP6oQhuOiG8ZwPaDCU8tIPrPRGSNTjWjVAzPRssbSatrCr
AIboTi2U76WDMiCTnV1iPbG3xjHA3Bx45ZyFGON5AlqiWicYmo+7SpkLXXOpE5lxCCIZIf88R5rR
YFPxV/4RHO/EocttTc+VxCe7a1amx1Y+t89sPBQ3Kx72xlJAwR7HQ1aPs+EXjO2DmcQX7wqw1ITW
VuN49A/WxbuzgAd9BBKZPYvxGic8PZP95uQotlJWJOz/nlrWRhGEs8qweWvXgJuRiWzTG5OdxBhD
F1LUgk9SK41meDfvUQsVdWq8DsiZDRzUYDwgwhtDbMeTQKr+00J+kKmapcd/RZ1KNYcyNd4kxhZU
KE9FfBr6ATXYSqrt2KxXnF1q5FExDmYrcGnnmWImrdQIj9Yu1b/jFbJMF8GDQGYSGHmHEATc07As
tZXvaiv+d4hfgrXzi8LbtllGMs0WIoH0rwU0RB5QsEXeJ7P2IYs9tS+1YqSRNB+nwQsqH0XE346N
7TtzHOAkXA7xPhYolsf0FEuhM9kSOqchbjWMw38Z6mncKLQLpvYMnGtwSoDgcOw6dZfrcthpV+GV
XGvllvLtkyvUZa+9LRzwqdu0RsLuVjg/MyIEhXpF4fT2fkDCazeU+WnjqiUzVc4o5VDZFTDKldDm
DDFEHokBlYRcJv2oXimrgRtC2xrjNIuxVtIcrA/H9ys07dkaXkz2g3c2JxBzscB70hgXeiz7ZrjL
iv70imsPu3ciK3zmsCu/ybo8Dgyl+JCOLCgY/eS2kz+JuMKaEalZ8u3jIQ9QLoT6/U73nx2x+P16
hnrNEqiVy1Uj01UxOhHC+yYewX7+I3kzdVhQJJog4nq6X/JhRUpqvPKQKfS/e6VxJHwKLNqMUBHE
s1eYgE92P1NtiSMhLs7H9/DhjOJ3kTw4441EKhBm3Fw/d7GS1ATCfj7MApbpDlUfxn3Db99OBSxi
UXiJOPZge002L+fJNulzu8ODw0dK5RyC5anWSES+Lg4RwbdBByE/crpDBghsppih4DuIXCNBw2JT
Dt4xL4tMcLQISPwPEpxo5mULEFiAWIqrJ1+DmUJbvYWfA5oDB8R1fe03BkyIYtOzJlf8Ru6uh0jb
n0QGSpsE77PgT5TeaGdl0QOkw3qgiabCEoWWPBGzKw75Fq3t28VxZaxRTM9nHWoxCWIUsq9GVh09
ABWWkFoRahkLOMq6WU1NWzje92tV/VPXCFK/X6wbaeFnYJpIt+eI3OdSPRklKZNskSnlY2VgKA8w
GHbfW3vRjgzdiiUCHN7FkZXfSMgeNrzqMi4uhrwD4urFwtjoZBVqlYD/UfES/Oz9VvL65rV7GTPt
96GSJaup8fyFqgz4AmhJotk7rDHYIJKM/x9olScimG0Fg7lafO8SwIDr3QAFMpo6susU0RckzTUr
cRSPHPIzLFOHzCxoNdRrr2QUHcxxUivfkPS+PUxdEo/X8eny5idUm1CmkQpOTeVEhn1o1tI1AjWs
WLsFhrPKj5YfhZbEZfuKpHupIKHuzuOnlTeKPteuXwMmhCLWq/P7tJ/Idv5C/NZIcYaB/VUOYeVP
/DESrjW1buEFKCxISkWEM45Y5WrVHMwaal9MxFmBbuUyqB1m1+le5EKU9NTIzYZ9T2O+U4sBdljG
1XUU4V1nUu1nlRuGbUXH4TAglEQt3EaYVGsjId/wmWEwi13rr3EFx1PCFAy8iQOagEvOWZlDNIKu
zcbnrUAhB1eugjqP1lSwqbA1rsJkdWmEfi3iBBBxsgWxtWEoSqzSV+1rtZRX+FMcN+sT0jLracET
833Ve0kOiiqXri6vq8sYr5p1oatZxgR6n1ilPbUdVdD12CVjjOXqUCDc2HqM+KCCvNBKipTb7b2i
9bCw10G3BFf/EqFW9sPwfhJIvfe8BcTkguowHRDnEzZWduvfhHc7EPHtjDWzUrQaQfggW3OghWAT
TPb7vqvHKzc5gQOt/72tvSIykoAVURf1thpzWxNb6d9lf2b00nzZW+UPCBTOezBhKQpPQNwCq8w2
NX/pUYrqXP6MTRkiIAEWBKdw/aNVRpdK0mWE/BdQqJ+zZsDC6TaksHU1xAgPHXtjjRjKwBQG6X0I
AKn9xzfkOhfgsd30y6aVCFBu23ydRGeYYJ9z1coUmIEVhsokydd89R0Ij2tYMl/iBzkMse4qPnmC
9GQp+56dd7X3v8B9qVPibY4V1k6Lv1dFK5r6b9NPErkd+SpV5j7SN4Fdh6fYNOfGlGmPGSiwLrV+
mcrcPknAC16jFmlduR0r5FG6IW4zVEY9Rmcr45pTfwpv9tISb02alvNKpWNOwh7wNBoK4IyCS7K1
qlkbCNUX6IU/2cLfzRRbtTlIUxUkZ+XJbhCxmK0hXrWOytrU3QuX1X3SrlOk8yfNq6fLW/jMTXeb
qjRbDyOtS4IPxy+xIiqavZ68nW7SEOE29AvyBnB5+qMirUAgktqKBQX7EMo9XR+bV9xOuZD1CZw+
841XoOG+aelqkzcziYDfxV75gao62/8LACLPahQI1s/9rh1Ir+/e3Mfn2hJ7Pi/lPdFFEi3w1Smm
QazTMvVab4VVCIXmJVAqBLl7OhGbsmPd+5y56TsXZxflPELDeNplYOskfGfT6PZRaJ8CItBEy8fq
31gVWicp1drFd3JR5qLZ725rwAHSrBAYNMf1Ad3z8o9be5FDt3YmzCUCeiJOvtmnrVOpCP3EuhUy
Fb1RHZZzR6gPy9XrqMXgKg8O3VB08mSHCLGHnIXljA4+nkEeZhNRr7HtTiLnKR3B8vzol6cRTyUX
o7E/9yS9kkeQCRhYZHnXRshxhgekBtoerLzPsETuoC3XeP4Dal5IyskRW3HRzuXvetg1M0cPy+Mf
UFXnY/smAllJiVlBhrZQJkz41d8dLVf9bDPsRVRSHVQeO+DOjTQDH1zolvZ1mNF7UkjPPrsL1ihR
JDJrnkWzjeYBamTSK4yKFLjTh4TWCZFwmAcvsY5zr5lI5WzHpVACkitDpDbx1+4TuvCedcNTCvkb
Pejci/Sf42tA4XpIBPwEnmmm7GLzbvrvKOWqXcD9rAwOpzHgaY4ZA5dGeklCTAqe5aSAoteFu/wh
PuKQEfNjMXm+CJb8juzPiiTXcezecvOE70zvGXM4sX/6iLqNLSRzY1lJgyvjzp5Jklk2NRCiWd7K
lmdHz5xAQW3Wtv+XZ2gCWZiWtkDVuFWxuPCTCewTZBD3w26s44BPaK5qsl1rAcHU1+WAmjVyRVAR
bMv3scd+QaSrrPt6yb5ZgLpEfMhSMDECqaSpq95WEuq1TcF2vOSvbVRxbpcy+j2kELUNu/8ZCKgC
1U6O9V1IOZbIOGd0aHgICtCPKmA4Rw8ywa7jldde13pf/LfA35N2Nt97uMWnSXhdF2O0bEcx/LzK
+7fOHiiLHsTjNjJyhIyrJWbL0eXmIMlkNCLJsqXH9dSplxkiyijvA+oAwdSR/6OrxzGDUf01JbEt
CzLpekd6LR7mNQ45xhW2I/xF9c32nTd9dHInD5c6h3drdt+r330SBGephKHVBsJIemJ6/tpbVSmy
JwsZUtbdK7JwF/tNPc4tGsHAU7Jk6mKrPoqtJOFu2SLypOt0AxxJh8Dkvn2JRJop9t/bITumDzkx
Dk4JZKcxzVE1cT9baa2u8LKIUTvkrHYJkiOd34VzoDftta1qBr+oyjbFme0Jvl7oMmyEMF9yHovK
SYlf4srp1IkYFdK9ZlmhM74YZIgpVkftK+3w8vpBvNXcYNg7ftQTHcuUIMlgzjojnkOE/2+nXCZg
62IiqbU67DQhE/WPqFUnH8xX+5xyqESGNyVCqO0LOUTanJowC/vycdOqu2EUZHGNU+iTEOr+nzzn
SPLkctEjqU3tKOZpt4hS06+90ZehQecE3cah9518XyovRSdAb+/mczA4L2hjO5ZJFciyP8afWTLt
rSwaQhw1WpXJgTsjYFTQMa8H+OjLKwLQ9MSGjUtK6d1EfCFgUNAuO20Wxp9lIxqNOSdahCFyRLly
NV4tC9Ul+v6yJs9v1uegJ81jd3yKBHIGoArOX024c0DyLFbszP15p87IxCXBfQnNVycQQeTGXjHq
unl7/Kavy/UOf+2ysCU9sk4MuiXz6cZpeao1jfoSuSHfBESmt1+t0YfgbEr+Ccyi66KBFVT/Bu64
v2vgZksnP/XGwko47IkisGfN4tjvRHxNjc8b1BtB66Oj2F4DHtR30g9JIX5+JqoxF1lGv8S8f4jm
NxNnNLi9PN17jFkr8K/lCxoEnixUEazA9TfSEUdCdIxa3257owkXysz7SzBAuatgREyRTPQPEoEA
4SfZJ2Hd6GuIaEd5OsCIJwyuOc8Ye9SZQT8cjf3upDI427oCQTh8yMZdgprSOnBo9ssKJ78l1flq
KIMYqmuEIkjrlmPamQx750QBKY1knvOGPJlP7KoJbLzFkDifx3Dd8vPKzAN3N9xMm1BZwGKFhoEX
shVt1W03ctVD4sWG7Kr7q8GC3iNd2yXMV6e7P7eOjfvEByNCTJGBtfud689gwupGLQfQ5dyXbEig
F6BikavLuFSz9c/XO8FPuplDgreADThscCkSi5ndu9fJx57eOValpFKFaJ7//588v6sgCW+Dcc/s
w0YsuLnBJ7a0ceCvx0Lq0FiKq5HvyLUkttlV4oIVIb6V0diaYAxPcUq1Z0v5Z6dzoIJTMwsnzsdn
93xbtKnw5SfkkhLEnjfAbFiXe5PWm9Cv0s6No5rbEwylXur+2XeakiPz0AzLfChl3pnINpKxK7WQ
VrzGelbBZfY5fUACPsRghhOqoIWuLblGSMiH0DdtA/fQhUICqVDDV6ZY+29UXyGpqeKSinEls+wW
mXSbs7VA/Ud4Yb3lhdcRQbWTzx58VvZG83T58oMayo/RRaqgVX0LXjlUdgAc1LRXhG7nsrrDYRcO
4yMOgaAdphsBkVwo8c6cPKBpc2h6NtWzisvrGZ7DANClPvYloJ5XVFlypzxXj5Xf4y7XKVAkxnB4
3+EQ6cPsNwE2QsErNM/A01vzQd8Tf365JovsFb/3ox2d4YoUxYqXXUcyV7ViQGU/LvjPnirqd3Tx
5uxi9GhHLbciMcrBVxY3B82XAOTo8CzewcbfimaE8PcBQRQin20a8CZdQ35/30fn6j+ErIq4YsOy
memIikk0LlEMptnN0/CTrlSLMBR7xD8NIjgXb76EMGrhWtH1weO2eOT789j+D0IICMD5TjOL+/1z
h2a4b+dW3OlmZ1LSM+4nKuHgrDpnFtA19x/mLS183E5SAbFbGtiw2hTD+ZI/FCt+QaMEEgMTMwEf
39Eh+AoDbhhWSCPzOlmm7iHJITSv/sHFIviWHJ3qG8y37Hd1ChS/fF2qLVGcEtNvBUVFGakPvZdM
gq37PhQ54kdbyVJto+V4wFzs+cu2jlLn+GtizWYMEBqNWW4+aRF8wBKak33kbDF3i+4r4C/OMzOn
77meb0+Yqd8GAqBmgBFUC/Mf5AklRbwi6s2N/fVYW4JomnAfLgpc4wcn7D0PnV9YFcqRIp04QCTN
ULa/ZoztOjH6jDFRp41y0KtcAMjva/CfQa+bpPwyi3zDI/2fSlwl959rsM8h2tiNG8DgAM2SUe1B
Lo+oo0Nhsi1QSWzPSzPMHIRbOeVnRjSXN0Eg/b5E3Mhg8dbMDhh27UbgrMWGlwDbzTUI5EQrLsxF
5eetAbgG/mv5nVK+d97Qa0m8Ii+caIF7kyeSDDcHEqKMeWJqZUWQY6uQmB2WXt8ojs6nzO9jUywc
QGUdbLqtlVgmUX7j9NxvPib3YpELYYDQGprDR9XMgvkdDJAUfzW/jzSYgWxi9pb11MxrO+hndJ5u
Z5NzsD68H+8Rs56mQNHC6Lmv39F5zSmglwIZfqkL4w+9GxIBy2tXiXunnAFwlhgK0GAjPX6uns3c
UUSypX4U/ayqLZFglJayovymLc0TT0CaL3rTsWa503CNciusuAiab9E1esS3Hs+SVkCzNJ7XZ29t
3H4c3hX67X/w4uGR37vvZckPLWpuVotrt4X2UZ5OfH9TcXVZVL7fChkx4mRtN7HoqyzSE0OWFb/6
va2qTFs0b+9zq2BHqIXr4Ci+0e49ADWhId3itmtD25cRcbCH0I/1hlbk6HM3x8C3lvPmBUgMnL7Y
1e4K0eSsPzecokHX3i9L9NvzidPSDtn+TUKZ8NyPrM8SmU/B2YmbzskiNiETVB9mP9bkQLMy9A4T
yLCJ1huhAnBFkOw4LKpT4QV1OHBXuP9E9fuqMknEGUhwxjegYlK/tWY1WvrGMIzAQrHtbK37ujMr
OdMHZJ12zctp9+vng+VJeUukL5oVXBYM/W3a0bQeBbzypkRCmLxcQKXg+16CQeASDTeaDxBbDfNC
v+F7OuSz1zdK2qsDfBuwwyQmZvk/XIfGp6TS2rWsoEt2s6UmPytmOSLsmf4Qfv3b1lWz1AZLCO1d
J1h8UjRgHKUAgz0zJ/PDOzQIGHs4NLs0QwPRazwb/loI5BpJzme8eVH8oY3x/0cwtI1JKPSxHL+Q
mFPMP26uTO0oGJzpmaEKhdfGgJyLWx6QTxS+6YqlyeGB66TYGGZbqldMwsPZk4gwgtUqvGki8Mlw
prxpdBwRsbBJ6a+iFYnBth25Rk8iTJsJV7MpOyNv68j+9U97MOABM9THkB+gfWUU5+9vUOtf7b3u
NYXIbxGI5FI2rgBejMQbflQsc9P3I/BLbpmmaSPS794sILUcqEAvMKUwxzZdONdn3p3BUhbHevYE
uzhwVQX/wA6PMOKOJWwYmuXAKnUw92eNDfFAeiyz5znyzK5PAxHv6z2/cr5YmojHwO4iS4tFJJ3m
meYM3t1jrX7GDVqBSPKOcnfzHDXKjI3F92OBU04CxJ6SOO2xmSIs00V7u/6TvGd049nAe8uKQLlj
6wxys63sqkfARsWZb9SJ48U4MQs/gICGSxacm1q1KaNoe+8FbV5graY0dGIO8vXReEYoNaze61Lw
VBf2KxH3Qw1Dof2/yniQAPGus8vRE9jDQmunumC98V8xOZ7yyrAtElomPloqeimyrr5JNjJqA2dc
VeKOSE8jEeisL2X4tgBBQQwSMWeb+cEh6mB66J2TRZIy+UMZI8JRUTrYqTNUBd8SOdmCHLEnx8Jo
jTXosAGCOx0G9yI+Lin0xklZnFEyD5+7rTN8xAC9Jx9DH8oNmuOgL7jg/JubxjxQb0ynzta6zgaw
qrXj59kfst0UyBgV0sBdrsMeL/IoKkZuqy9y3goxIasRVZ5+yLv7otXs6oSzfxBqrEVPPpOuNISG
j0ieXaF6GgybipMAGq//KHTInuHIri53CFvnVwPAEF8BdXp5zIC0Mh10sUnHllX4BOXqynbF+cbH
hrYqvexd8U1hD4iQYkFm2TDn5z4Y/Equ3V505AyPza6Ct/I+GJWR3e6NH1g9AnT6bKUykCLKPhY8
0Jw9PgpT3/GhN2dxB+oWZiVAXv6zC5I1DrTTpEmlye2x+mPFHGEp8htytX5jHZcfbZOKg60d+xt8
XPHJrV4GZ8Fbgb6qmFzAVfvayBed1/UJxIWGyVyq7HeUB8lPxlNTkKZOtCXLEc/RG/Z23z4RkRvX
pzbKrBrXO31q2BeS+et6CY9t3L934oNDBhKO9C8TtghG0nTtkfaOCxOTVoCZgjy09+2/KZZyCEu+
EahSq/GeR0o1z3Dl7ib6iqWCfPX9Hc8VH4dmgaEKyMEqQu0r4z+PFNL0W6e8ejoJeIfNIPugeImR
Npf1cUtSvLCaEjO1OGOIxtOzOPMH7Gw+e1T/TfqmMAtlTtBtSykQASbQXV/94Zk74DNTAx645S0g
YszQtbPxvaldzNQzO0c8qctTTfJgz+kymSbWECZ99yoA7QYATKrTNbpmN/1GlCUIlRdsGk0/tDL0
2LHXPVYYYjspQzuERKoHN5lMJHhMmpPKw4VW9lIf5hHeUOZxMDTsmnTec40S8s37FWfO3E4IkLd3
iAUzBMMRiNPPd1xzZgYPMN5Kk+6A/mdaj/WVwm8mjCZ79QQUVushH/3dr+Ep0mNhpE/RLGqkjZJ2
sfwLFhoXBO6dAB3g+oJPvBYO4wUGhkjZSl74tpo1Xl5bgS7WKMkMdI8eN4yn+frJZo//I9YhQBFa
ZroD/RT8nsI5Dcu0/mV55/t8U5/MOKwHWrtqaKQ38cIUWhxynyyytfdR9vK8c8/1CZg6nT7iza8o
AZDSklNdjo52Zo+wGaLINKUGkEehsj6/7trZT1LF7nZhkxObiuOlsm07bV3eI72M/cMNkv2YzmI7
If5OvFNtDVDyVcdEWqSk6ctW9tWbVNrxoOp79BfXRWboqRLkfNpCNZcP0z2hIITRjpSsmIocMjTK
7a1wEqsnR06VZsZPnlIY2owCxZzhOVzMvt6OfCPeiGSPT+05X55nbPIegdKlHlGwYC3GrUqv0fwc
NzvZ6DPD/sbV9S9H8HN4cxo2aRDTWKJsAVwFhT4+4ntxsITdtcnZsNDH6ABqtNW+BKmjYieEpfRt
+AqUQob+9x9Anae04OxZoPkU5JfomYyx1KGOfMU+WI3P8clUiPyTlznex/FG+sdUw6TtcFPOMHc7
qxuYTzFOSF2uHrJpuPmCB9f/RsuZVdNjHNo8ErL5YmrN+TmLYH5PtP5Ktb03gWs5zw9KfDtpjw/T
pUUx0pzXCjlei1dr1I7rK9Tucwl9jhuFX9VmLKfpjZiiOVrqzEi+09YEwWJx4XebVA3m0JSnqLP5
cix8i9Detm6QROOljippuG0+qMWB0n7mEv7X6UXPi7feiGEqrNYcSI4XKO7I8kXBQ8pHvN5pAvLi
VlZ5tdNCjX9K+L6crd/h9Ry1tUuJftHL8CHTQkXf73Zk6IPYrfE17umQYOf+aB+tvD0steVZUFoD
wuc3/r604EabljNWaV9WmoBDYMHZkqBWSaPTR21IvN0BMM4Jd0n/y+Jc7TMOGrAebR0jE87kGZkL
P6AhDGkE4LSTZiSWLzBhzXMtx7SUUmX93WOHQqEONPIWuprdwRPasSMtWAojgAgnZdGNCVrLWctk
ONNRrJOIG/udrPO5iA8a2Y0E4gIEH7EEx8t0E2nRfaWul+0M2gRlZwAAcWsn1lequhjgFCNz5C1o
4Ci7WlK11hmt+cLJ0tQMIIkVpFG0bv0XadZjUZ4+b+ccYO+pFs/fJgOFdA3hjaKSxDsmi18La9Th
NcC8NPAmALPl8zoyDU8WTiJVe40Bo32Wc1Kp9dyGNX1Eh6Fb+8JUawbFhVvVf/wr20h2gDy645lV
ewF1yu+ffbQOfCgLT99BATFhIgLc3L6EJ0uK/k2eK9sqZp1cDWo7HCKcfxZaCeIFRQ8TXjjEa74q
r49Z83eKWiUhohDrSovkbs2khg0oniVH6tVWRqaSoS52+xJmAKE1otujqGYJn7FI0k7uo5wy0nxA
z9VdgY4K7ju3bS/cgtJHtMd9BcnJjIsb5aPDl1PdJiOi7DssTts6cSIdnwv2QhbvO5okFQN3AE+I
8nTfbmW1Ddvoni8wcRyO1n/sKCfHGO3U1Yg07hs//2nVqz1FfdDsT4PV/nvuJXwaSEMJXkDJZxXD
0L1X74hC9tGj0KmsvMvGkBddakAGBP2sZp8uHHUGj8BsGD2SKJePnMfZDnq/nUmRzM1w2vQlw6kl
TnovrYPoPHU8TTcV/rRHYBWJAdTZiUNaqfCiBIzBpSbYkDuTzHkEHZ8GQ/On38aHZWyuBWdcBdLG
e2TmoIgxlUMKI2UaxYHVQ3btRmfF4+2nqEACHTtTaUnpZiQz6k2W3IAwyXqK78LnB7J1d0Cue1Yt
r/bFM5vD4o5TTbbu4XFM9GQaIsdGGm/f/dG8WxscrkZIZgtqTq2+4GujffJ9lwPwvVMcwbDDLB/S
7Uu/33XVM5PXvOnJOix2dY1KmDiUAkHAlxhtmPVWFRcTlfQtTu4VoL4ZEvYeyLRxKz/bJo4GbXtE
zEejnh4CRTMyWa8hyPORoJrQmpb+5y6nkj6XMyo4Uahibvsri8ALEQDiGODIbBHWNEZ5VEGtP+Xf
jTvs7h+bjRGGaR5wEkRZptoGo7+jVvYuIcLqcJKN/5+gXP2H8+ws1risN5N5aKuhH+DRzi6WQgzo
X8QZTMx9tzpaoszkHLIBmB/QHLdbCV/rK9O8xtbwJX5ZypWMG7jW7ukih3T9L2WdWlfKCWHjR0u0
33WgX09T41mKvCwaEc93fX03dwWWAguXBoI8yQlGAQsxEAAHqdx79jNLZOivIZ+ABDHMn4g6OrTG
rjKyhPRXH/iOQFupXSMaRV78z4Kw0swHkOWXvcuC+Hq0ruKclhLjWK5jxe3rIMSt/amRTR/lxDyy
7G7yj+AODEQ7mHzCE02AdqaAX9RDVX5EBJX9KDJVoSuCvCus5Mek+dPf+ayZ9YAja1107nMv6j/D
WPa1jT0Mux/amvVDaBVzhLj+E96NW51EnvoqCtvAaxKDkKZeI5ge1Ov/OfNuGyDilcoPBth6EqG+
2s2bVCrpDcvIBDbtuKnGiw13rsq3gWzXVj1XcCeQu4I7sohO7ak3bo6aOqL+4T9mNUcuPkq+hu6y
c2u8v8dgczfIOmwdxxBH5n2zWW+D0ZzZ6FnV56JZg0ntnsYWg2+sz7rIMs11kOw31KiU+y32nCFL
5SSmdKetORmUXO9aMk2XfRDjXrZoVhZ+326VvpRpXHN5ccz6HRi5I8sDrs5jQMscWnKyti1rXa0t
7NsGwkm5O3GtYeF5BP+pY7jbHH6mrg9i+pRS7sfd7NTZVQgKptN2EN+OVl4azlWeTUYJP1uC/Dml
MwU0FjwBOQKuGbPw8ElJ+POZd6FEECLB6hruO42CcbkKZitu6tv1QEMOUHyj8obd8J8V5qiZGVRH
t3uW+rH3xDTZkojqh85FF1uwykc358TVqCFgSkFhYid7SLpSdOQOb+/vY2IB5PijComQKqCGN8md
TpEc+MTm2myjlkTjS59rEiiV63PIeFt4EjFjSHDLkStJ2ah68Lc7H37hwEl4RMRpcPRgsbjQ701V
H3h45TCXTEmut49RLWKRHczQs3UtpP5zOEJSNJavHVPSHI+BAuvvdTkM/PEaVjR2y+MM+RiHjj/V
DcJkC7S38JAtIoEmKxIwSYSPOL5yINFlzF2ZTwxROFmjJDHgjTtIkMbk7/vlrhve/Ei3P0IlAZap
mJ0w3igM6ELBX2aQqEyWEpmrCqTdL1wDY1TVA+A6I5gILX6noRc/NQO8qBxwrkk6EEqm2UJdORfk
s2UZ3wKUxrFzNYNAK/NjRVDna7qwJYjsc3IF1itt9VKRKhSS55MVdJP0/KYw7umQkQwplHPYEeu8
sFs+6mEIw1cdsZqWmYwTA0kzJk9JYRFmL4VHZX2b2AncI4Ox41QkCoMNazH6pkvk+ZXTC0fjbmeD
lhz4fvk0ymiGaciwOqw1Mk/ueCt4KQWbQbneLG6bLRLcce92faDWy4U/rtKn0jmhrkp86v6Addna
tI9cYE1VUGiN9NlWuih+opf55y/JinYlFjB6h7uxQPDFqyJfxlgfXpJ9cAJr098vzq8LY9LtXDCl
5NZtSKLkelHQk/3QtTX9W7WxKS53KK3yZtr9EzsfYBUosh8pXx8O++EV/Y1b71cMzACtpFpVzt5v
VSbYhx2VFkh0OOtrzt4qDjktEJpmsyaX9BogFZT0EqOPTR5joU2jdHpmPjMzaaVsiKCqeFzxHleb
f1EOWu7uEc6fwqwtIUq6Naw/w2V6ilMYLyv4NIGwFpj5TpmV6Te2pcwyL0bGGyuFInYWAaA64ewK
oan3M90YvUYUjroIbHBBKLxMOixrZktj9OK158FGTLaf2xmu5KmZlMeVCpBegF8nS9LON6aJNPDB
b8UTgByFMe8+lg7NlnE0OY7vFAP8PfhDqonPFBXhi1SnGIQ2nWQD/jq+WM/E7iRmEIRgXBL1y4kn
EWdgS+k27F7HHx5usY2rNeF+pQMEe1DKhDeN6tpXMiYPWKE8JhmJCqJHfUFOUjyJAmbMvq2uib9h
ZXfQiGFxrsrTLm2fIgMEhV3f20/uJX+a23VQxrBEsxIHgt9bojiza3/c99BevnFxwkZQLdwTtTh+
mt9D/BmVPC9zeftnfq9Er+fUicp6lXZy5LxDcYtCvPHksmnFW/wuuYkKfzbNrsraBd3+XiDWtZTq
EX2cEQE0IuEttC3vNDaDTlQji/1eKNchEQmSGNcBzI3xv0NbElflUqI0RDICZI/KHepF6feM5ee6
VogepBQ+RL0/UzJxD8nr0Nt8JaIjy9jo+JAEMr7tgOAWorPyFdTEaRqr9VtJvtg9hkPS0HDUBjCZ
753+i+DnHEHBPyVK5hVa9MWJB1fvTKsf7iQEqVBlWDBK97q4LJI9sEbWdodFMH6SG9G1oV230Fmg
QVLoxKD1+21EcPjWA0E8HvOD6H9Q0h1bZArjF/88jfQU9hjCmajqmG9H9yxoJCuVT412aCRDKLma
Pcultr1xuuOthCwYyV/ary1VwrwWEvkfmeP/mhps8oPkUhmgT7T3yny0aA7bPuoXZpDgE+SUhqxY
JJGYrcFOnldps2Boy/JK5Mp8/ea4MkZTmZto4DGmf5EiTNuchvOB+2mLgPv55Ey4sKRtRVlMz3nl
OXyEZvpsbseT81E7dL759tKT84rFy9+M09koY2uOMApAXv2LbNAnZpsgHDfDUaNGY/kFYaIn8Ssw
YbLv0QpM8mFSkC+MHZDREsUG6AZw2Frs4IdOY6V1ijLSC5M7NActhrIsGpadPzVws+pVXV6qDIw7
edAjY/5KhNC6DVfHRzL8Szu1F6HTi36GHEBv2BR5b2s7/wqX2TWXeF/cc8dSfPOMO3oALQo2cY2e
UuY/h2cdjK5/1QWnksQMAnnMHJVVAQHadg80zJiWsjA9Rklc2/ucvFN8GhX9D9Kz3SGIcF2FCWUF
2RB1l1pZ95YjNjyGfaXQuvNCH0PQf7HMKuJWO0tt8Di6cZGgMEMREdf4ncr7ikuDluHzH7vcZuMQ
UuoAfANPE+pNK1wHUdMTTPJqnEN+uB0iFpMo8CWX3xHmA79N/XQ5xHAjfFyZ+2HyGOi1l9t/ytGq
ZmhEpvYejlHCacrbJAA5obnzJBRl5DYsnxgbwsuUiTfaZfCy0+U/VZgIp+eTlEkVjmiVLbUYb/lQ
xcIKz0detZKsop2up+YbnF+5oo2Yk0RYCQO56fXsDaoVo3389G3j/cMYyKtmlbei2qGGQBG93UFr
kf2DMnREYSXadVFc+O52SDOce69Ul+wq5+0Ved1yKqVj2IqTF4Pzwzh1etjv/UYuJ6RijPx16g2U
FKRofRuiXLvQbR5HPVHt7/RR42+nNF/c3z5mHlJqtIlzL49+thw8kC6hfkCVfIPjhVNbGG2nj3t/
/argAHDzPE1051GFS2bRnZHZsBhQPwfpK6vxDZv88y0GVuk48aBduo+J/TmoMPoqIzJqPdoiS5a9
h+dSBKKNYIG9YK4UISpg8KV5KVZVuPzAz0SPVDWB6mOWow2kdF/TpSlkxHpayFFPC3FK1BsEVeyg
lRYjQ1NdxfN7sFC2E6orwh2m9HL9ckV6n1GnEof26Kblt+MlvEwpQ/n2HbBkbzA79Oc2WPNl4FtW
G41H7/2nQ9S/m9jR107uurhqA2WCzVxphy/8t3kaB0Ep1XgAwMjfmkrVacRI6DlyxxWxBfCOo/3Z
NVZcSceBQaXfkq0XpnyKqrJhoak4e+TivaoZGx16Wm+IYtu/K6G6z+xkzqyg5eXRuJJNp2pu7mDZ
wMgyWDgiDS1sG9zBstMkWM+N0mnQHtEjOiCFQe5eYFVBO2q2qCLZIGeCHBrCkZGIC17Gm4BzpkOG
uFV2k87wVuC4ghHRuXczOmKY4j+RvDEXBd73OfXHm0mJ1HTBPcLt5Qgicu4neEmMZ1CZdaez9E3b
+A27+nhI8Kt8DcvQ7hoVrLwfJ4siN0GYOJDGC7rwJZ/922iA9y2phB78DszzTPA0gVjUqw7zDGzC
MZXWY32TzFXncj6coySHOhMC2eBHgLEg/M5ltFyof+8GClwmvA62BwFvJaAvrzuEsRX1yRk5uIeZ
Khl396QSm7TfX3MNa3acR/Qpxph7r2sMJ73+ZsLibrzNxivjHd77Ls2YxpNuGbkJ9FR0ZWjB5YZP
rWd71vc36/IC5EqU1GkDb7ZjysQU6iAxGWJRG29/JaWYhM+l+fC6KzzB2Qaj3o+DTQdzpCOBXZcQ
F/7qIUyxiTxtgVjHjqVPddf0lthqWT3SBavHY78rSEVJAMXAo9aqI/WghzjCLE4Op/s8OpOOceIt
8E/315u0qC064cZaJIF2C1bxO9olYA/8wH7X4DjPvdyuhS7ZqhIRwoKTH+P48FuRLcgoHWeA5c+G
ZvLTyWKtmA670WiMKU4bcrKUUZeKCHh1XE4ovGzRkEWVlH0gex9+sC4sr/6jS5Jp/IyzOom+0QYy
La/mjDIUMxzRAADcsNcS1wd9CpT80Gv95NSInz8dXH4bt/1UFTu+OeQbSU0nlh504PoEX+aHAui+
1N4Ye1nsw6erf3fvNpi1QLxhPtS81oPnbNvhq07kf65m9x1JkqXdYF4FQItmTpyNDwnhONeCqH4d
Z34N0l7txRt3HEc1rVujyEtVYW0ZYRFkkpY5F9KhBAC0lp0iIMiPtIF+Tnt5fHDnPH6yqoDtsDmM
pfHGcAFY/0xtWuM3IA6LHTG960svgntDfM+Y3ZlJP2365twPgzzr8W4HR8ubCVeJwqEdLD0KeXSq
3Gq9+zdtmEvXWwKPUGxGXE5zK1xuGDPMz1pSl4xRB1igoGTLMOAUlqXFwGi2tNBpKXQyTrlzTd7X
9FSNqNRzCvAdKpXuWnd1wNTaRBIcQrFcc4KRjWAOBqX4pH1mpr30Kq1hzAB+dR2XHeLanoFf2HBM
qUssuZMCu6CeauKYDTBLSb83GjjS/CSuijtvB+Ca0KcKwKBMTsT8EOk+LhgrawBPZB+bW5e1Y1OD
sl3o/zDHalRlzSoEibypUTQwgLWq01GC6JdwFNqs6e6PyK7OiuLPyGgFQM7zJcnBmmP1s/qbWZdg
Lwf17VuEM5Zr/Pb8yYFhTkWfXLm0GtwvucDnJ+gxDMoB5D655i56dU1Spy/NMM5STaMo7/U+l0ny
Rt748vq2NhY9kreZWiOKHct/oPptmsSb3A68oXc3EZSp4WiG03JQjTeUhpH6BekIaj+R+StPKIvE
CNnF1EB4RMq76MEKnWgE3/a8sqBEf2VCotcsaSYZUG3hcYj5vtwY5zGWNkiG6EoAkyK4mTAblu11
eQMl8niXCc71SIdQg3rOC5NFNU6xWOnT7xDvgYjV4MeUQ9R6Jz5He69tqBNs8Knpmx/otYo0ZBwe
JjJYgGdjwJsUJKQUJfuLd7jlHYN91Dr6SHHb/Yhpiyv6J9KAaDrsQEgeC7pgyIGXvSJjMxYOrxuH
ySi8TcYT+vvp82NWqMwtfPmmOAvcaubMO1WkvDQE7RBnb9vI9SGtbvcEriXXykPGdVOAZvyfmdho
COgm3PnHyDMUhPsI0MBWYe666TvUOQUFFpB1vAvcRQZarmoLWDW+Mg0NpipV6MnzyPYoNvTWcJ4r
b1XrJ3ieer54LDHj/SEnCXw9o/rlIsstGDNrHsjGpowurKe/ts/0ob113W9fLrZKSBqfyXZsl3Cy
D3eoLNcI7nl3pXngUpM4+X39vebqW7VAZP/6/HYn6xetAB9x8wr5JSoHmm4g76+2gmzWgPKNP3Mh
O0TDnrfySxxJr/1C596Ke1XqbdWz/clkMykZbPPb9WhGMFtAxSDJPLqERkKckVLnXcVL6k0SMvz9
TB2pdpYUIdyU3ToxFFytfLK+epulV8Q8x+amUlplmcjaxvnu3agpnk7J6qzOx2Yfi1Rgi7pl+R4c
mEiJ6HL2LqslNUm9w/rfApqK2MhLMnF4RkDECx8xdIH+ZZ3JfGBdwvz7Agc930i32200mlFgAVxq
0xpYrdmujrw1UZog+/kncobzc0SAsTO1Tl+N13SiEsOgyKykNiV17vrfyFb76+uQr96YyLGCSa3W
ybpOqkHAObRQFfQAv/j74SDwFNT/PkEVamn98OZ2yel4pxf0mxa+QgisYSJf5dVERHVeFWBpzdyT
gKPQVuIdj8pm56xMrc1VJamcZ98W68lS174dQFI/ZWltRye2CrlLiXZrL6YNetw8r6DyqYosNYyS
AOBBhEUK9LdP6d8SNPhTYOv/xp5h3T05rL3ERp1d/dN9EtRpQPpCULIXI1RHndrxi6dEYOLAa5RI
tUXAwASkD6ucyCymyngcfgyjmBFMIRzHzvLVOzg2LTf+kFw+QXMCvLOpStdFvV3hdT0M0R84XYWN
LDeiKRODuTz0aMkeAf6/vbSVEnlxZ97StwiJAiVeM7HM5famOga3kO7JrIHAM1PHiTS1mm1CmrW/
wfrX3e7WoIbaSO0QI/TBU5Su1JAsM3MAHLhCu43PuI2KZfDPGFwda/nsRW5RlMFUVcsbS2QsA0uX
3qybPECquUvIggGQA5aBLcJruBR8/d158JWhOK8PqoCMTq6+hlcB+ed29bM7A3PGSQpMswlNgAo9
0VIlZdtMbsuIs350IN6a704nGFErCvsfe/v/5ejyUTo5Wj1dgqlvj0GCoqTXLgH0p1/munPnFsGL
RuIt+7s4iNpomeWOdPWMbSsOT5kE/zpyaVXcGDDJUpn65K6Pqwhmu+zB3JCAWqDXaaEeoZnt7TpP
uuoM2TuMIIhnUffrwYrjIZeSJiZ4n04UGTzg4MYlaswdX6TPpbAbRjhwwTxpEyIujajC+/Zxify0
Pi8ewkmnwZcTzoiVLZc1H1QGlko+n8nFyoIoOmhMSvZTJotLvx9k+NmPzkyATptPL3siBC8loSGq
NwBrV65OsXSdVloSdIUI4KTK99nJqlHRBtr/oICOBObxSUw83MnCA9g1bgGF1GrUJipxGk49POU3
o75W6N45HwBGDSwu4TnmfZ8uBeFr6kk5kFnkPZzL5T5GlOBeD9944yLLzYsPp1M15Bg1oQEd7y+m
z8n7D5M/L0aj4V2/s4rDAD3ANURhjcCDxaKHxZgqw3fpNCwhIeXN+W0pk+pmdOAOk9BNWDNkeUq5
i+tPk3wmycTvz9iJ7jOMMomYOsXIDC7dghJNH9GPlUnqbFaJRu4AMCtzpWn+j0IfCwk7s1Dw12LN
yhQlF6fBABJx/4yyM3qBYNTzLYDBv58VbJLhi/sPP+ez6NtM6oLGV0GkWhLKp1LtpDusS1/SAinB
OWlo1m4B5CjJCb6wVfQTg1dO3slon+tGAlZUi7ZoI5GITKtrdUzUcoM5Jt0dniy6lB7owB8w/TIm
i7B1djbgGCRfNYxGhy7xuBoBFYD/OjG0I09b831jd7B0tUj4sraFeuSp/rQyumqcbtm03P10e1IG
DTVAj96OBS3SyITAfKXiSC7i5yXAZxl1LaKC3LtP2WlDNjLPNAJpD6bxCo88iB/RyW/zSkounooq
yh+NcXTTsZp/6PlDXZTV1gJ3pC0PRPabF9p5siHrnxl9F/0lrmUV2NtI0jJObuPFvKKYTBg3XDTR
ZGI5eUi2Ik/HLlHocLjIdNJhOOB97woTj3AD3VhDPtuI9SThuiiLrkGPjA96lV8UafdSZwSTPS+J
6KZmCb0ThYbgUaTf1gtWiZNvsVpPVKzoLhSceI4P8JAr99U1rNK26V8JGtgEuF/0yWJj1PH1BPfR
3ftlxeQfd2/x6H8q2yi2Z3yGMmDvkVibqglHeHfLKYgLi8eVEl+w3VQJOM79Oddt4bMS9i4DTVfR
TglPReL3GBAp0dGWgsZnv+a9cINj4PfcbeeOTBQAFDbXVrF7+zaqbs2DMhP9EjVQU/fPpy0TGkzN
gdJUvoYjwwpBbX21Yfd+UR0Oot8QziJSb1nZLNpdmHycSyY5UAxy00eQsAcsHXUvP1JSyswfcorf
JQyqqMJuX2Mb89ybML9rwyHww01m+1iTXptpIGevJg9GL2adoJ+MShQQOcopxbOeGpdMKTwiYotj
GgGXsCPsnJJrXxhm7X/BZVSd1rOgolV5T1m8t2Ypx0ToI+IULSQid0+8I1OeRxDheMgz8FSs8dZW
pkR7OQvYiLz6Wp2ExH9hRavyRnM1g3DcQ1aSbDPCFny7+2ixC4d0qaVGka8eTeF2+Rzn8o9D/nTW
djDOeItirXrE7ophFz4NLHG566XP+lDWzvUPLLg/fV3QWUIc1IKyVBd+lMgNlvQLv7FQAhPza/EX
5oJWnSu1AvLj/N1wvN2Zbbyv0vVgTYINMDATt1GhJHw7wgxNF7wJeK3vJxEKhAQflfwZ+Wsw+h6C
SKqakq6d/MeyBbqWPrrRfuNPxPNJz1p/NnOHqLi9atbJOc3SfdmR4ucXho7KncF1MFJ437nXzDZy
Hgwphd1YbJAlcgyvk/TiP9TuDTqGoO4UF5neM81fOJoPlgNS2sPr1NXHeUlnob6W0AGiqQOY3KGn
xL/kUxgH2TFp4EuqUl9KakuMCLp82gIM1BvDAm86aUHpHF1bv4CCj8jjAfM70ozownGtHI1ICluA
EontZabUG4VTkFHiQpFsOBdY6bRU2aynGtpDIJ1UjC+Fi04KEGR63QxyzxJ9YmrjCmq1sH/k89Ej
/iCwf8tpnpOo6oP+okXDlw7wfkKz4KIXw5Bnn9tV8b6Lf65XqxMLxmyxRj5EcowHNCypcpdc7SVI
9ekznnsWvFflg8vNnfcyoFJD3k0RTHIBnDFqRjKwbEvWxNyF9tH5FTuaZYovE2+9ry5TICxzepw7
CzHVJDbA/0RQxn1lFKdYftxlTQBLDpUS8JVXLit2TVeQVntZ5rrkF1F0dpiIUGrJYVYujYNJ01rm
NqtB04vMs5YI3oQRxXMe3qZZgm6HPmnV9tKvaQcG+IzUZkxvbjHF7n8G6OoWs+IhZBXzx2TmAtGv
3Wwb9hsZLHGNRn3BDFSGMy5Id18CBgnqXDcRWNJEZMaQVO3iSXka2BbuENBF6MzaKFTnWry2UwIv
bdmCmCs6u1cNeniNV+biSLcvYlDLA5umwtUQ35vRGZ+DnqKPCSZ2ScYnI7TPcw/Qnc2TU2SU2uRm
oeVWiMKAQuxRgTsikHp8e2gP31mENwzHgTizVVsJxVFhL0NDdp7O2bkRDm/+A15usoeJRbTu0HIl
a9lpUXWVW/zsAw20yoydYAy4u/vQ2HBCERerA3HbJEgXSEOyiTV7XSX3Sam9XuYxuzx4VmeUfva8
66YGgHTJNMRK3osbCqLhjAKYCSkKnnHQSlsL+oViRNwbg/lS1P84qAXBcGb/1vsYDWHcDkmV3BCn
KZ8xW/Zar8HcDXAFvSBAOZjCO/JbLUj1e19CUkGnKl9LLPr7bxo1dP3cV1hPUooT/oTmxyTGBLkR
vwIhVTBz0A+T83gzBTQSSjvKT7bqmFNIuE/C148pvIXYzjarDrGDurFE6flhBrG/WkcyvGT072I2
DpbwIx+8IDjKBbcMmFbbjvmZV8FIttxGAv8m4ZJEYvZJviwnksUKYVUMOfc1cVOCpFBiC3Zs3Cnf
6jH7Hry7HcAL7r2+dBtQjHiC/QGZ1QdW1uCNG1XDWRr1iDp5JJFurL7t10RdLUPkep/4JEvHeGz9
QgR+pPjNWKCwnEmWwmAkpRDs3Bp8lQW3DFT7UeIhhSEYkqmf3olXuj+y9QpOnI3bP648p6Y3dVbY
ox1Y3KW8jUcWi5ay0uZtPAsiuOU5FmpJdJv80OghUL1TGsipcUIg0NMU0cAdNiDvlNu192vyq5rI
nB67Q3jSCEv7zG1zYNTwK/icSI5o81usTHjmlXA0YtDdg9V+x3bOR2CFYqgmfSiDPR2mQapDEEyg
D8cZrfKnDbz46/BMa38lbG49dkML83N160MgCfQfiNAbUee4WFr+L67hq5Q50pNToX3IdF7UeH5m
DHOcuMmybALRRiAgX25tMqDRvDW9Z7qWxyIQncnU2qn3mAV9pVZCVhpCDHlJJamPvHayDpI5/QMz
w+xOYKAsChaz0BlicvXP7D+tiGj0xQUJPTIn0ELLjTTxpqYnrYj43LwuHd/L2OHXa6eWYnVl8VKx
HB03MCwUpyZIf/xZ6oiYAA55p9Dm2EIA6id3HySCN21dc5elTFK9vwCMMU0kv2XY50Tv8YAuVBnI
JSGUFv6io5s5lQR61JK8VJ3lZ0RzhdPS4cqD7K42/K8niZWxVprkZdjZ0u9Ee/wr+xWPBxNeGA9X
oY4RJeLY68GC4WsmnOhb+KHtrxmj2Ke6ToWeHJDQVntXw3uqEo5trBKDTyjfGfl9CN7nQRtwcKfQ
pArewiQzH7DpMhihagGMicxUInnJ9D+EglAy66qZWI0Wgmv5B19v20qUgATBLqGkcG6oIOzk47Lk
Qf03hXvQJ5JwzoxI5HOR3UKkcDNWS+xYxJLfA0PwKF3IMgVgER4UWN1LuFziOSPJEznrULFdtIP+
9H6i1Lo6d1vQ1+pe0HOKkxapY7+rm+IKydu2+WxQ5PRFdCL0Q/akyejS9evaEc8TMjGIn2Wt0CNh
6HEfnQBt8/aXCaDiqO7iVU/CF/Qo+aiV1GeTFRHXgGQ840VBEpIaH+UScqHTUfSNo+kKWD9947+5
WxmW11/CF40ABHpQ9wmr0WpCnuJAssfkkGlsdJCRdvFTc9fQfZiTvKX/xkwLkB2F8PRmeq9w7vSX
2BxGGBFHcofjt1gjbIXlRJ9zJ0VLYtIyAzRn7uu6d7qybQ9vHgsoNjyogodG4U4TRlt5OowLAFFD
kHUMfHs1TGmaEMWs2U5qoBeAc0vybRQgLwkeYvvcyeIm3DZCEFPudLEjxXvig9GYaFz1t4UUwZCX
DLFRJTW8wY018rxU5woeUC8snDBlz5jzt+pnAkZ+kLmHq3m/mchQ3TsTvYUUZgJZ4d/VX0Jkry0v
wutcRAgDH4pYXNYiXOhDDPXFHH/8FI/b80KL/dBJkeTZ8HunrgggvtY297LusOdvZyGhRuJ1oMeq
U3p/rjcyhDKoD6TOlffmivj/li2AQMYc2UKAiMQvPQo85MZJfEP9+P7n+q8eOWPD17HYHTU/CL1d
evWQChEYJ8WPZXMXydMCZaENC3fMxqmnImKU5E/CgUuj2tLGs23mIBDwJIbES4DFUR0p8OtuNgcT
+h/fplYcLzPWWNWr0DSeg65oCN9iscWE2CoZ8MZw+nxsnluKoTwmfHJhQQzlVxwBxSK7wMA+A6O2
aAaKOCpkHFDTkAopRbIf1vV5+MV8wZaLaDTFeP6fLB7OOlj/zj7fpJ3Bo7H462E8/76qKuLvXaA1
nB/CkvXlJs3Fz4q0x6Xg0wAbaMc82XbVxfoMOtHe8hgj4ThWlT7p0OI1Q4DBU4mqDWT/WqEJXKQH
6eXF3rBjo9sDpVYRmKcKgMeKF7N3UZtRwACwwUE997AuYobCXwQAgr5RpTKy6KRCqeeO+/Gz6wRA
TMjJGsbyOVGaEx49NoIUMgUYpONG+qKZkUqHRM5Gv9r1I92YozOuiR/ldJY0rwfY76P41ugIirIk
y9o/rVDjlfEUNlSNbVl8aCuVlY2nqHeSxaHoTXH/o1Od/aD1BizPuZlVax9RZhLYXGtVo6EN43bX
VJOExF5dOvcL6E8nb+9XBj0v1k+c93ECQUTYO/we3EdKanXA1Py4VxSj4u7BRbDUmu8Of6we4lQ2
SqcdYr5xooyn5Aq8nyIVlRjViEN/E2jK1KqNHbIu64YJifSHQKdbIHDiFGoRL9h/Q0TbCBk63UVl
kxgkU6gcSLFZGeDvBYcMOy9EUa9VrUCsZfw1fOCkhqpQIbqtXX8ZH6jkGF4lIAkjkPnrBqj2dyYr
5NFPjRJS5amoirBtNtVloNYtSif/ZYKFDJsEkqbH72U/LV3+sAsxQQ49FNX0mY9LsdcO8YFUVlXw
dE2miTCiomBIDC+ODONQYUkQOJYWWAYBC1+BSz4men8ApwTz2a44wdl8S7Rrr3k3JNpT3QpgYYjI
Xrzgwc6SI21z+IIMrIQnbTKKjrk39v4AAlG9p1Ec8Q7fLbtzv1tGhdEh5bs7sL5f6dLdcQw3bNuK
e6BCOfCmgPUoZSmakQvaSdzMDFrRI/HhHHnp42MD9NssAfY7vTJwNzdZf+71eeeauL+sB/oJ8xJ2
adKTr0Tfq0JR4YqQpGddV6ZP1u/arTx7Cjb9jwvEZrVacpfy6pnvi+/0B3Ri2CsM8MRAhx1dPlKb
xhaQRB9GjaFIf8ftbLFKa3x9O8JclvmWBccxBJtzjz1kWotfd6KRg/jIgIqqT7eyilEuhL1TU+Ic
PeT2zzzzD2Lhz3V51I8OCjB8DVmO+72YBPI2pyvO8jMQo7gaJ3OLeZBbA2gWN4P7BP/Ph5xutFg8
YoEKmrRBWTN7MGL+Sitmght/5n7q1GmTnUX1Y4WA9x2/WsFDJSVBHQzMAJHx6/PzsvRGuLy1YLC3
tZUM/Tz+pjxnPN+jc6DQRQ0spVBc6HP6OunfJWn9Nsiix61um8cSaKTfn5zrzPXvL+vobwBJgKMW
TnJUwCWLFwOxC64+/bnFAog6ebnUODECteTfpc1KAEnGHjGRgYLtF8wD4rgsXjQhBBXklcY+i3hJ
ZQUjHDyK+459289Y7c2/BfZ1/EW1GJPhiXIIfJqolkfL1KomUIV5p539IyP7H03r68DUAkXa+GJd
1gVjOsYevvaSGnHdCSMH+uhw4nmzsixpCD6CyC6iMsZbXBE8S/7/spLeGWqaNjxb7yhGJa9qYLAr
o1H/6VRE1dfoXZVEis395PaWV/h1nNcaD8L/53FB/8dWl/6bcVkfcPuynHQIDFl0MRb+F7x8wyqp
gduUr/UDPI5D1aplIJTJYkcPpMB5ilpvC3T6lN4o6ztVFiQLFqr+8isTV4jvsLL09/PlPyM7yerz
UWZ0IUTnQAPn8zRGp0xCgz9WfrYLUKZTCFLI8KRdXdYuiQc1HWohH34nkpshoDoBErp84JDXYWp+
jGUwEArnkvHgNqe4xpi2tZOCpVjlNJZzkCYEhabbPt1A+VQKsSUhy3m0B38X4Ev9IV3Kl/xa4vzg
D+OIF4A+PPdCbWmqHSx5GMbit+6B99Cgc73v03pBnb8V8VD0RwMHGHYZmeMxYSsPQ2TWD+/T6fsX
XZTtj8ZaPqEks3Lu876NOSjxDFDaGV6Dzo18p/H/rrF3wvtVhczwFdk6UteKT5mRkddnHun/ZJRC
oSvmBlrgPa0D2EpQ46S+VFtOFkwmFbf3MPuaTloLGsq2925hfRgh9+el0sgG137Hf1j1K+3h9Zfs
QT2LhMKCldladBnHnyodIA3lT7cOl8TLVQuSBNDybgqTHevpC9Wz582Q4N8u4t1NwsYzizhxTTmb
Qof74IiaEobbbReiD2WyLmruP1jb82rAfDL//gNWYVcQFEsP8OhaooImI7q49oHZRTSrr+M8/4U6
j3Dx4JyE70C+kiYgP/NhTRm/YGNud/oebzQpCQkooICZOJqnoOO/WE9wgUk4rJ4WD3ESNhStw7K1
RAyf2bi7JW1Bb5Z1gQ62KtkzMmBnVlip8Rx8C6FxVbczYEp2VNsTZqzE4Hwz6mlubMDKCek5jtuC
sXknFv7+CvrOKVKe2YekAkW1WzlJ+KyvW0oIX1weWE7ElPIEhWlFron4Z1eFOcTMXndtsjggaGzZ
GMLyLzilsd7AvYcOvYhQCwECb4u1NZ+GyKscVT1G4E3ckB4kpcHKWLaPFGui3VdwozaZ93/cmCYQ
Cu12+IlJZZjb3ZTKXgyk2wVQ0Ou+yG6f8eXLw9bnksl5ZO5cEoRR7tWbXvKleEriktWxvX2omL3/
0XiT8LEttp6wLeTLk/lWPTch9aaPDxPqdyhhnh6+J5N6H96Cc7MUFX0R8ZZim9LjwsyubbR2NO+J
yzVkVzBv7hjZhP7mYcOSiRJifaJWHHHKYRGtNer95XB1ZnM4f8seBdtanbLpIXOAs2GeBJSF/G3p
8Jw6JUwt20Je16YkzeFJTxw+HfcJzBsQjaG+l1jLRGDIO4VDbTdvg+RFSJv9aMhgKxsrRMgK3K0e
b/ivycwx+Vlng1z/7wmspoOklayKEq0dn+bJQ/Nj2fv/HXJ6y1MmGt4VqnkFxTxJB/zaS9W0gqAx
+jCeMXx2B6FfG3KVZi2XG4ULGa2/r2hIHAqrTKl1NA2WGzibwfAyoy8XmngqNjP1/CynHQ1FUZ/M
4gvmWP7vi973+6+2K0kbaJpaKRqrZeQt3FTcKOz4WpshwXbjgqO+XTYuyrvhWybWVMbXenFQVoFO
6KNhaUKn5qNwqkHnQhqduKK3dS5TgosADo2ZQyl6kM5asgeg2XmIZRI+KJ94zrMQy7H0nbrvMwil
wa3My1gTVK2pJBt5y8a42PJHvOLCLtIK62XodFCo+iRhj1+b2OzmpaBihX5HsirxwUdpT2YWLraP
/buapt9k1FZ/BRk+tdkMpoDV6yhGan7EUYO1k58W3a90K4U2UC5tARII0iXZhr3eoUXLPUTH8pAd
XJv3ylhWIRGUNtaFEA58SA6/+kyR3HzJaHPri+iyhTetrlLNoitqAtdMmoJYSnhvJU+XLq7N54zg
n9Ne5B0S9UsgNJme6CDrB4q4CNBksyetiZ2Y2ht3k4DaimiSURbrF2uYTXY6svNIpzWQObBnZaoV
NUrQ8Y+rA3kNUS/U71WE/YL4ryvYsmfPJV2F352n+P/udFvdk1JiUkG/dvG9veAaA3RfZwhusZ7I
CLesg9oqHbQiJB1lwuvVdMVpyfr5hqhJl0PUWxMIKmnJRqA0Aym7kR9ecp5leHf47rcXOGoZ6U+1
/T1WRq0lmviUgqPgvg33LHW/tNo/6sriGY6PJqz7aOZ1NwlD0vungnzxsnwiCqq+hej03m8nel4g
TY3T1g4GtwyBkWatmcGtLItNNq55ppnoGXgc1T9CIH51DV7UK403mSys2H3/lC8uXYzXteoVv3wK
4n2o4CnCMZBjmJP+Jv6GyDO8RfNcBRfKTNilisnpM0BQ0ydXp6LLIK+oESgJQpKdcb2duM04PDSo
IROrm8x/B/HXEfv/HbI9vakmQMSLCvQ2DueWmwHhSUR1ylaqOXxwAg8k7PVp143+AwMFw0h4uxi7
Eo2RVdU7yogvpzvSRBxFjo0IpAlTmjjxArbbNVsvPBpq445wf9CEq61cDRfh3EXAjXWGei9iD3wR
6XEuseuaClZySA7+bciuw+je0XF1CBCFV9sW5lYd9EicaYj6+4k7dbrKTpswSju6NINJ4aXRHjyl
jzcD8BfZjp7gLcMQ68tCi8rnN9mlvwC/1vyRnVXBy4Y6nfdBot0LmsSJQW8ViSVvJdgQEHdypMbT
Lb9poZhqxYVF1ynYPqCSb70t6LJyQosQL/+9Twa23gHa1ajYGvrqw0sv4gGGmOEEQF/8LJ3xYiHi
H7QVDCJWZpK0DAPzBqxQ07lD3YVIwmV3emHR58Xp+eU3MvMs5aiUqKJgXdIwYjl68TKep87HG7ZR
qvmnjxou1DFKjflAPpizx1qKFVn/HP3EStsVg/ALDTC4nbUMS49y0dux7M62W5WlKTk06Rpj/dB4
iqwBeWEUIHO/rKZxIQwlVwwch6UytrOavZS6kEK/lW+9wO2Mpj4GDTMm4BxZoi3i8LuxcIDfkLf8
wz/4XOuEFobikTMjihvjnyo8DVuApD6dWd8EHwHxA986dgZpd+bx6eXtHadIx/TLmlnYETNZGtC8
R/wXXwIYPXLuNWEBp8j0ZE+LTpdbaQYV0dz96aVYe2x6Nv2hQPhqrCqRhzECSprE9uqF4zlraO+B
b5pjPQheaeQJFxPhOnO/LBJ6oIesSupiNhWUiMAgwx5lqUcudlSabuSfj16DTakcjc4+G0j8suKa
R8OMozNUg1xwwkdCPXe7EnRh4bPQOdKmYeFwCcpNa+vyFSqXuFMmO4Bg9cCLmEHqRMLjGkn33WdT
/alGM9TYaFYhl2jOpViZ9IS9bX4teNkI6lM/zOseKnJ6Qw2T/FdoVkJ1IbWplwHvpARnB/JpQF2b
TKo2em8+rErKh7sSwrbyGiYY/jQTmjKOqwgEDV1jeXtedJlbH/cAQy2buO1Aqli6zhas9K7wUEoZ
26sXV6YfrkMcd66fal7E2wRSquGtMf72QPCovdykFHHGIPbeUqvNlc3BzA+nCxMIp0poZPsrSJ4q
JMwIEoSL6NJ1S5l25kFAkerVKaqIepRSdeIHP+fH1UaZxBX2WDlwod7P57eNJ5HWN9BMrYXDXF5e
ET+kP3uX+gfH42nI8Wa9xAcaWWbmvXMPwJfL1AqOR1XSVbU691CoLnePV3blhw9WdvvIAeeTYfmi
lXVXcwRb3tJtRaDZDlHvWcCjYU/WPfy5+BRVf4yMWHMf2MDLlVg37+dtOiG8l/VbdT3daBKOt5kH
/iSDgxMN6t0GN7fKQ3mEppjfplmGs9w8/dNDQQfMUssfYhrs9isX51egjVT5wlWI4LICNuOd48M+
WQMiJY4gHxCW7QKF55BlKAx55aWPcjCCG+I1NeNWOKgMURBvhXdaKhuGYl1fhRoAkQQt7kXqrPw2
fe7waCHZT3+yEsXTqLh1yGZtwtj7Zv/v+NYfbNzwIOh/aK/K2EVCVe7ZuSLG/GYQM/OIWiszlDPF
FOftNvdlDCnn4kh2KAyGnjUGACO6K/vA+Q9IDbv50r8mJcH2gm0OwFbCKENXRrwOewmJ3+45xjkR
ehbpYvYMw0kstaMNgetUJzkUBdsYKHN+hTur+KZivsmJOxmTW3wI7nI8HjEgfT5Wo7Fe+3TBr/O9
gQ1E2UD/Tv5SfXSKquBux8sdVqZ29P6uknht+EL7B/s1sWR4N/1xdBVx7wZy5EdnfrA4qAdnnYPQ
br4NhoAUXjIhvA7BAGo4XL0JmnNFWCkYsSZSStpvAnJU2fgTIjYLpM25wonAIYVKmJaPKcAqZXA4
P5u3WaJpBDfvplCPZ9TqiULHSd6lQ3+J3U1yUKJSNuOvKvMrba/xeeFzK5FJMkDX3qWQI+qcRoIf
gCVK4tmTPyV2XOq8kFJQbmD/1bW/EInErH+40S7kMVqXviM59SCHoSLz3X6LLYXParypGcS1Q1Nk
OsfYxkMoSB8rvm2kbE6Tc/TpqRokUoaW/TdomdBCUI0YOfauD8gOGLUwbjgPGpMSrGwh/G+XBhVs
Qsp57I3i5qX2Y3tR0HFMDqwqlMRsj7mVnz65BkUhHCt+i7tucCMfMpzdy7TWAHDExWHjQtHA7Viq
2ezH9TCG0a5EE35BQBe6sL7PJsdVhsPbpP+gN8SiUDU1si6tZMaDncZfYnXPQRx3FvgpD59Yjv2D
unTd+iMjLfvnOliIRdJR0PYLo1K7kii/JdmstgKRlzu6FtBAoNZeBi7r7646IgmiR9yhvneyrTXW
nm7IOoiHOe9ebGYEt7ZXYu4rlb10rSpkzku5jKhhTYCnWUaOJH/VXVGtRaSGZVCNrcU3PWf9UJEl
WJxB6HWBjkO9FgvJvads4ezEOW641OSVHZ/x43EE/Z1xxNvLzyTY6gLNoTPWl+/LbblgbDxA9ij2
0NXuTWRvCPHu/sZrPmZAJAqARJc42FgqOvHQadRSdPO4IFmt+SC7+xePmhowXkna8TgUlH4gWSaq
29WoZCjLePTXF1h3TLED4TVw2lofld0ToTDIG3HZ8TQh6k0rIRAuylNk9b2jSSVFzHKKOxtBZd7u
u+7sbB70IaSXX3DpZ5OyoLQ6W46BJgee2ve+/TdqA6lZGuPG9Ro7i9sE+w3Uv0sOlZbXoYHD6RwX
tzcCT1JoDHUAAy3xUmHImU+bK/R8TCQOkXJagT+bmF2MroXY3eJYYuzLwIY4FKAif8w8ERF03E3c
zeJ7OXmFSnMQ7VQnZ29oViFnAl9oHfJBekhFv6LcDEusFHWVvMK0TNtc5ZGXIe9Mcx/VRf7EC3it
PL7RfgRHi8XhQOGJKVxqUydWyFV/J29BDaWtIs/6z4w9NN4mOIwsvtBv0xUBgls6sOsB9dJJH5pH
DB/KCVWb1Ftg7QsNNT3vkKEENZpD6/+rodF9GTYBhoAREjXdUcaDGtohKSU5l0sUk0TGm8fxKmQ+
wRWZi8yTegsqvEKSNa11MqtF/dcC/WAQMHnnwfDxvbwpYzwuTCvsMYCZZxu+IcY0JnFbgsYdQOt9
2vW4YtDX415VBSY7xd335HjJghlj7oCDLKct2KPd6SYOs3/UPYs1yKQkpLX0MB7TXyvunKeyZ58u
ViFMeW1r5cYaKgfIhMFNE/y81En81Y7RSMPhhWTVF0txK3bnH1TNyc4yVMC2DXdyCIt2kYgLU+Gu
BE83HYaCXve6wRE880gPfyo/knKPCSvaacfjGxE3pohp0cOiOhwIbrPA5MSjXwZp/s3v3eI1S/LS
KkkKjEYl0RFKuosd3kZOv4JtgwYYaUHtOFSiIJsGyyi3frpPCEjqILawWz23LTjZ5rMo+1UFSRc0
i6s6+Exk1TefhUbjL2Pz353BZtTzesDt/Wqxv78whpKXNUlIggHzDSW3cNzFRpI+VrZ05lW9i1TG
DIMlaLNg9d5LLpO5Z8ctru9zJeJ4u3hqxz3bKMgSpe4Jscpl7rWy+Wp60OfD6VrtRIuZQ0YV8GbW
g3GoVoYtxJkXx943HGT/vj6dt9GV9K7+sIrvKzEzaeff0iBRzu0KrbYkbnIQrMHBdBCAPjDWbQEC
QOdSFQ/d3a27yEClAeEo6Mf0QCkJnOihBSVyw9SZzgvmtlCAP2ycQx1m3gzkC6VxdnEuOp4+E2Mf
dyA1BmwEKgTTu8lRVeycGKo8EESadlA15te5awo58t+FOklAgKxaSWi1OyuxM25Zl/zL3Qy3Vmxe
skfpp0Pb/M/fJ0OexEvHvfBQFkMnDFuRiWZaKNKqUN4q8XvAeAMnXd65HD1lZfN9EYWxLppFxJph
+vQLMw1MW2UzxuvXfdP15axa/urmQb6dm6bPdTKpwu9bPGG3TsAG2ds8XRg47pKyXO4BCVTZmuvv
ZvA5gJpv06cBRKYAru0IdFEW1GBaECrFQn3bk+um4ZCMcaGabo5fAempySKN5VvSbPdYYJI9Vder
ITTu/2SlWNwJwbW/o7AsboHMfvsAr53f/5s1naUv5eirIEl5JhU7cjO0qY42c+e+fACc+1LLNmRz
qcIGpNyZgDRyL6zErpj9fdWSzsN3rWcC9wqXFkd7T7OpIZBuGprS1k1p5bnGVAVUg7islBGGNeC2
GnkFMvu+DjDydz+YuhSy27cjWKWTPk5FUAsH7ITi7GNglXclsUclnAbegLePCkMtYVHgjq89OY8d
uggyzmVS+Sko6mB5EdXBBxKGG1FGvRkKUYS9xrT+m5vDtxICUAizLWAW1CJwPuozBPyXo6oGEQsZ
q6vdoezeuCgxZn/TcCnXPaL28y7RlMd/ISeSG+Z0hGR3skmetwWfOsBB/j56L4Ze6OV79beoBoyC
Fxu0oaA86DxEK15RdUOYiiRitj3JoY56SyHxOoNCCxCDQSIFu77tUozSuHHlXpZqSCvfxOt7Dv6F
XAD/4msoX1wB0Z5wcSUNQ9TV94gqcycZiEqwY+U6uPN5IC3+3kDBBnKqctLmaKLu4tTkw78C+27R
WToIzpf3u0endlTQ/L1IhvIcKX1AYedAZGeaYyzpv4kLWgppwhSCtgJKS6vzpHqbzR5vkG0UnLqw
lxsoZneUwPV77apmKeEEdj38yOtnNdGEGW+RgyRWLWawJ3wl/A6QW1DcLSjeYNa9Z9asQfoSRjRf
2fGVZvnRvf34DewhQgAB64Dv8lb+5QrgqLF5R67gM/o8bUacUMmrNnIRPgCuEcJCMr4BEs+/nmLQ
qrpTYQesVuoC0hcVDr2ECl4GNZLIPGJm5jElA9t/szmAKfkwpSZTKYQFCDoy/yhqqtJ13UexrBmP
HcDiMnzsHTevU6e8zICeb/rk8fXL5ZZiZgtMg7gGxdvgRl4LqZwn/Mx9+wOo47X3gtPDHnP95NfX
pkcZPNzgEaAPBWb5Ok8AoWr8OvpHzLgQoXD1heoamc+td7PCahZorPRc0i01I/64TG67z5g0HY/V
Sl/1uqafuOR1YztgaXtSppDhSb4FZ/OIWiOmWArhWCRB2ViZbMrRAnQqvIYrS60VINEXEAoEN8sO
YgjRl/NMBZdsN/XMFXtkx13XVjgT4H+1z7W9YREJCb61AGYDg8zhzhAX9TOF4HTcjy3nw34LOQ+/
jyR1ygneOm1tRO2uk9VY00K+1uN/BQBgKjYTolqwY/px6ITI+Eypj8gAZxV9c5WbB8If2Y/Ne47Q
F0LhrfauHoLDXYuG0+8AQJreJhVvbYhMRU5rFXCEAWEuKa24bPF6+cWGYBf9bGQdXF3c2D5uVY65
zslnLj+LAXTVJ2JQyP0eY3q1HVnMFiX1T2DVofz7KySFbJp3uyVesRMOZPl36neI0u6pWuXhtzvQ
uWWOr0640LV9mqmbCXM92ROF/DydFIqY4kVl8OP2O27Feu0ZGezqx2FJa4h/ZlEsDqQMCmGu9bz7
KnX/77jYBLO11ECEQEkPPVOquQnt8gp9edXRpiOg/rRGVvB35uli1aIh8qx854t8KthaI9X7ax/t
Mpj0ShTtZd+3Md7+5GzDyslPXoTiPhZzoETNsJ8tta3MtcKgpflJV1vEFNE6zPMxqzWG7CADahjd
98PWBTwUcyye2ZVUFZygn23uAJrgth6VfhmFIjQJ5azWKd9VfxZMHb5bs4SHyDUuhApYV2TqkXOP
gVoUWqUX3NMeirJD+jYTNv6fEHau1GCmpenIKbSi+qqF9ngFp92PhRvYj3QYSTCiVBan8qOKSqIB
FzRURWZJV2EvfWRhsH4uo6qrc+d3OcZ7UYLdKQwvDKOfC2/zXY7+VxB4lVEneBt3463dQmgtnykx
eK85WRxYl0OZgJu/4Xm+w+yqpzCt6dodf8rl237M6VaEghJbaKQZHhNulImc5xUlv/DHj/N1YqWv
o5lFWtYO32YARV7N1nd8EB+KpN/LE4TEX0dXFIL5tEnmYq3vxsQ9rezFKBTVF9gz+pBfYJ8oHz4a
V7fBM8ouRr75cXfpuR2Zz+QiKYT5/ZC8ZfMgvuYy2CbiK+slJGp5qkDcCTYhK8rxQpbSD/Ip/Htj
FUKWY4JC2W4vxfOSfn5JIhGxI6hTtIMxTD4A/p2tO2Bssb7qvVDqkcQR3L1R+lpRkRLMFAPJg8RZ
d/pjY3W2SXp5dKCYW4gxwf+/i4IQjcdjYfUN4YFsIsi6jQh5ddlRT3ItdN7qDuG416CnxKg/LDkA
uUC2/BQQgJ3s4hKZOvplmPJPQAUs7Z1cMhFPXmc86QcEdrc9zeMT7JUzVjwygnjwrgZoNCqx2IHU
E71JarGfmgNp5wlAV2TJCwYmMaJFvTsxecujgzsvcG0ei1BZL0zpws6HV+TNZxFKiP4dptSmSB37
owa2b6dyJvxFghIpKcfOKW2jo+VdDBkU4mIMwCPKsENZ/jBV2lqnKE58yW48gX6rIpzvfKI0np/X
vGTyiiJBjOrzvzumCH5Q7xgshGU8qPKeQ2g1o/HgeC5YK4RbC0y1Z+544oAfeGZelqEK1p3gIWIM
1MGDqd1gnSlNNKNXYiGXIZnbprrRnfSZO6k65A5WAIMVy1vqK3PiSIsgQdsqF2pALHbNMcRf+umo
sLT4poMwegQM7EZvlKIQnCQ0PxD1ByJgdZfA1z+LqoTfI/Z9m+xyc1dPhC6zGIAqP/qPRenhE1sY
Wdm/7zJZImBFINOyd6GHKuhqr2LBXuyg0+5eLd6rOR2kYGWSRmeWTxq/oqqZs2/xAB2JszYelfbv
MjSWaUDdJVuNbejI0fsFcBQ5aMnxVGQ/uRnjA6VIrTDPp1CC9XZ7x/kcyjo1mHN911w1VRGxSxI0
IEdxPRvkPjZ7vk9Ac1K4mX12eIvnhbr0lj2IEMP1TBgNDWOuPevWhdWyGYWB2nFFn2D9l1vnsmP0
nKr3yngi8tS+M5RSkgWny9PbxawEwVmqOwK+VbiTFwPvzae5SVpXGaG99URDY+Zla89z7xzYeSD1
23kC8rjqIHearttRGoOQ8ovtIuChdtxm9fyX903oE8eglfI+TeJA2d71uRR5jn3Y8FI0uWhkH+Gm
EHeuRQLQSey0gGeUkg8InGBDbWrT6YrO4nLyeK9bHY8EOUGCDBc0Ew06reXL4nvOI6FiW0xf7C8G
f6v8CoFe7/N5h3R1SvYLydpz0UQQ6GpuVUH8+XR4/V7/nSuJC/4qGioGQtvA7n6MyjWqVOB2ApmL
FB2Ov9tmKodXnsuWy+rRcOz1Lvn5eAYTK0i4R+0LdbmQUOeXCvdKHM0u/QpUy94n1Emht5yFkjz0
aWgSaUHbkLQ6wCnYB2F8o3PcM6ufySb9xs93bzyzc1O+Yf79PBiMzHR5iZ7VrOZ1tD5SYm8R3K0R
yLkARmXP0mtC19gJAZi0KlFXu/yYIaU5k2J667P08e2xCjsl2ky/mMCGtFSBcH5vy9Gv6F5b7xgf
1VkBoWNq6NzNz1tI964pCsMjj4zShFYWJpoqovg4SENX5lVLGL7SOczpcaanYU8lCW01xh6QRTyo
WXMqaAz70R6n519NhSR3Ba1ave8k3OXJoauP5pWkEi2LQ8dQUIcF/TtI+0/O2JoM6UitWM7LOud/
vo7JULKHu84y600otyEVsJNHnOknJ81vc3w8H9vvTYQ4Z15vl+Af9OKW9+bB/Kd2se0Vgr03r3oV
rsJs54l5nnn8opGJExzH+p71CXa/HxxvkI/sPAxkfoWOoa9i+d2UP/AF2iMzyRKFy6cJCvEaWfg7
232M2BIpQQZfKThN6rUMMWETQxGA104yN+WMcXdX/uCfgkracd/KSz78a1rkHQ7W4VCve5qWdkcS
TyWMR8+WjsxsFLoEsi+3nHd0nEMpvwnn1eFZSzS5OXWcRRyhkgvsgNKYIILZYFluPQ6LUkSzZ8MB
IIO628mzbXnWE7l7W8qxo3rN4bD3Y7H5BZDiln+4diggHdgqqM0csY4V6+0cwIzJ3Obkkl5KxEQP
h2PBU96OraRkUDpiQB5bAM4jUvBFPYMKBAHM7RGE2XU6eCUjVy16qJc8QfW3jadmlABnfcXROgXd
Zco/7nh5xDzTaiyjRZb+lpin1gJoVFrJQH92NDWN/EUOKZDCXW1IQdYP60nMS/7j6Dy3aO9jWfsT
GnK7jsmyHjotfdDancx7IqtL5EVXcyu2wkOu9Su8eGD/V08Ya771ygXKh9K0o7E9x7nphY2WrEqq
uggCRNx60jdZp4QgXMhfesqkA+ubadNw1UwogA5PYF0n9ulzJOZt3+/WuZ2+klGohOmUnqICKFG8
GcQTcgajA6nFDGgN9ezRLwjlY18zOJ9e7sMyw7vt0xcSauy1oIoTyvvXgCZPcVXhC/rz13zP1Owe
HhCrFi52kZbrz9WTgVxfhzFA8rrRNaBkF1l3aZ511bp1/TjUISwCcepBIhDDeHFm7jkIvXDb0yp/
H2Ry2lOaSzxAM4vtEvdFoPTEznkQASdR+Mt/+KOESlb+GWnIqVEOYbxeSinIjmYyjcPjpG+1Ti+u
oX6zEcJjsgwuhr98ib0JfEi5PiYw17zSi2s1fOUdExUvTyK9+mrKIsLDrYAGRp8VrAHvwin8EYgI
uiDTm/wBuyt9apGnpFOdFEci8KZ1Ot05uWq/HDtnZRYB+JP03Zo3ZtydtKedg80sTANAVOOKsKMg
HgS6wgFP/ObN55wOqlI+5zlLFoksehttH209PK0STg6qBjvxyvkTCZpZ/GCISxFiVpho7oMvfbal
1btlGYBBEuJjQqjayz9H49ObvBix4HI1udhHMwW+xTtH3NAZYtHNuNmfLQu4r4alq7xo3UYmb6AT
h2mzaNUyYfeSLx1g8n4b1XKNx74hiL0EHwvSpkGnRfiSYNC2uJ/w56Mr4F3qnwJLuvd1JtLtID5W
1FqM9VSS3hTlFWIPEEKT6sN7RvFAEQps2B6XsC4hlljg3Aga0yCiejX8GbEDeBBB1XS/H9FaVjAc
VxNy7auNDzWbx9VeVyAZgdoDIWdQ4rEPK8j5O1NISrUlWoPmKPvA8M+at9PdXxIR3DY0DE5KTfUZ
B0XHXUWBc4dwpUIUfqm9BlNH8xEjFMxkDWVaCxcLP8Si2szCui99r1M70HbsPZf2Gv/f2XJ/Bug2
yW2s+njK3Rc7s82cUDXzcK6YAlGR/pXNSBJxU8uxbBUh7/AeZYOvn0W/b4WmDDqaK69TEZOaEfzO
004zdNTmNV3hV8xB0k544WoBnSkNq2tkLwJLtseZPRA26zSvSx0ZcQWpl6qVl+mtco/WoBctwz2+
N9croyPB8QgooJTckrkfW8pVnIyg5JW5h6Yy+qotXcDwR1baNAci1qOjkP943YSjQi7OFjWzdi/g
VCoWTQqFd1Jl/9s/GDrwhxkBSFyiATDrFz+9qT1kCvBRf+BVIsRN+NVObQ0oN+KKfWGdXtI8e9A4
YLXWOt9qtvCCMsKzfpW/8dCz9AyuIgAmQ8XSDjbqMcSyuE2TdNsXu3AWV7oIRqqzB9lTllMmYg3d
IEIyhuDz309iK4FrTVBs6P9FAp/hSqwYpkI/BM94j1jinK2K5yXSvJ9FM8nWFXO15g12KV/QMbdC
wvmbLqWuHpUA8aTnde1BrwA0/DF8ipeNqh+BUwcOulkAL5RdS7VbSxAA+sCFE8P5fsa0fLBirCHT
Jf+gYU28DFtp9s4JcyA+IL+78rwq/XqLiv4IqjHiiGPhVk9da+M4lp0vXP/nVB+GzovXB9ow7GAE
/iRa+wzLPoRE9nTpKgFvYMp6+Z9eZaZhVAHyj1ktxUOSc30dYgJj7HncTVXGv2Ban8WWx6yR3BIe
jT9ZCbfmvJHd4tUfyLc34QMKSb8IEzAG7t9qb6u/u3zvZmlzbBUIXNSp6Tek1qtbxhLjtKfrTxS7
/AWd7CbLC74JDzZ7LLOWdsWcwoBKUJJFtGWt0M9pg5NBjnpQKum6YlWmvKcvTGIN3coLdSNyKHPS
H+Nj54CBNyGAs3KEnH33ZgngquecdlToHOkQYu+ahr1CORQucUq4n5aWLI05FabtiudbF43md6e4
kt79xzgdR6y5CRzxrpbi58PXCgOxlKhsN1qeyYuLMvP/IwY4oqoUlsKylsRNdUKWpp2pOcWAs9pt
luCNi/3h3vVvd0zTEiYWC1lWIMQbeRlppCBaUAiR/yUM4E8baHO0/gxASjQB2wl3pKDIJd45sDJD
ad0PooYCJLOWOPGFHLmgJuALobmooDESFxz3p5qkmZhAvija0IEQycmXG4BZH4IBdknXbKhm3tnh
v8/Ym4ry40RKi5pTxtxXtOtuMMTwvt8eDi1AhCMMqI/NJAa05XXO6IN6bVMXs1ksdTrQVTGIENTA
BiEwxjjKdI0cTMytMDvsCZeKtQa/hn6rFH0RhbIBLK8GABjWjnPsngkqGui0cWPhtxGF6vOnXLb1
kMKAqLInpIL6AkklgRTP/NCFdzCprgOSMe1/L5nOEondYiT+XrNeje2MxWxFGV2TI74CFb8UCRRF
W/TDyhW+GLPgJlGXXWnETsnj7z+FaPnJH7oy20zovNX6iDrA0CfciyqQzFqGw3HARfISetuCz85E
euaS6E0EpjRpQs/poKX2+Lg0BhI2raRxCKWXUV4lBz51NQ6bMYnAP8UrfArjRZMnD2jeWT0da2om
cFKO8qJPIADEH4StCz1p1CYkX0QCbG3TueHgFhb+Wt/Vh5tAtBOroa7WDGsotkj71FgXwaBWDuY4
hLDeMaULYB2Ytp7JFlZBnQrlcRs6mEPXU+ClapXreMbTdY0egqcJTqVXt2jMhQBotJOg563FEccV
SxIAqMHjaRZnelIxRnEPMg079avu8WXh0ySfQppE+z7TfBYNBiprDvcrdLhebway8gxnPPj1RRDR
UQ/FmdvDF1Cb53llEj3BlU7E5PcHOIi2yDZlODmQR07can7pkrpUEQPLYm9/xa5g8/fWuJ2vmW9E
Jl8KTPo5C8mIvAoD7QMQ/5+xgfRQ5R2gVVGPEBTCBrxsXOCMfbVHc/FxI1eudFVSR1U4UFtEcLal
tXNH3joxSZuUCQDGjEL6kW/Q+WpL7vSdNku2CuJqNCAi2hvmjKZ4Tgkg0ZGLJSH44b8eUGnesTIz
KpXN2w2j1IqEB1+Yle/j5KUg1j9je0ZZB9UcBnhGuF7MskLe1Xpn2Sm/2fM7OaIDF1WdhtEMj6aS
hmfWo9ZErsWkTwCv06RQXpVyNpqGlKdSN7OGYDPLaMIYLk5UzUga8vUeZ+u0Ao0WK+3ffXEtLplv
M8gfQZAVjATeqigZIDD2yMW7UMu3Uv8rgs8lceFj/fZjvreK6SWWboNmMDdYr5mT5lzu7dZd7+g9
G0Vo+g5l4AYLZjwS4IdS3rPeM7tBu/Z+bsao2+2O3iffCaMo5qDvFBfxAF4acQCHyeilONtkKlOd
PsWP674qm5Pa8n22uXG4Ifkh4/V9tQ/I1Gamc0UCK1pdQZf7DWP3lw/wiL/KgHlD5s/LahRteqh+
KQ6OdhnLPpRhSGkp6I+xsx1VNvU9CdjHhENcuEFJOi8hH3GG64bcARw2YNVFEetX7llozwdsqxbh
JO0E2uUz4HjVWrKQC1ttd3TsMANaKIZ0uoPawMuzavRV4G6F8h5nceoe5kKzNpkkBfwWKgJmQL+9
21aCI7j628IE8uBqI0mSc9IMzJjEM8E5MOiT/Ma67tW1duRBOLL7MoI0W8xPHEyFZ+6RYP7HzIXk
VeWdW8KWdp8A2DievdXlszx/Ul4l+aOorUUCuPnyGyZ1q3Rr1bIM1G1zLEIL9N8qC6dhDO2LsePP
YlL+q+76V1g6sW1+TGuN/VynHsYbkfJejmFJCiuEBjh1tR97J21oeM39STTe3WyeNeWnuhhGOZWA
TxvDdvXHi7EnCxfq4cwbyYIF4u8n5X0eulkcYIPTHcuZNkT3WXMMtZfZ7mTjOu2SNT2MDnckS65T
amtiwIVHOp/fnrr5InEIXKv+ms54fp7V7NZ84MDXYwMb18le9tspVEIDlY/jme7voY+0arl5NlUs
HhNyUwKxp2XoONfjQ9XcfUJRQTNfK4Nw2ateKSKSubjxjd3FLF/2aVzqopOx0W8nMk5+M7A1FYnI
ukPhzSIy+MsAcMgx9Wr/BG3JEk/WsdfCLvA080YX0ZS1ZeplJkwFbQ4G7rKpGKDM8nWUmw7KTZRM
K4vnxYbwy91sv9/VAWOFjmk4VDoyu01ExhlmcYXACGWNXW5XRrtH7+3fRvokrqzYdfjH/2/tyUhc
awJpaCDODGrQspl3ChfKm+F+8S5Jvej4B03ErKr4Ud7+u54Mszjwc5CfZ+2TKXUuPX1OulDwU5u+
w/4kVAA1JAuS94OyQTGplx7tAUOm+4m2PSDVyHbsMTar36fxcatH9nQr2OUsUsWF2Ai8tQJHjWAi
wpMCFJ017hOJq2j1k96Knnc/sTZJGgSbhXMcQ6hA3IylTsiuUbAdylMSudsYSVfsHg+kJK0+VsDm
90deFSWZwpaS/Lhc2WJUjp5c6cgqFWTwSsOf24SOlzWVSqU4FkQ1JzG3vqsFh+3gH5xYxFeZYR2K
JYYOmSn+wuGmbJyhw4n3RU6f4ZBwMHtonDaWXFjABOJtVHgy5RoSu+WQUd6PTt7+Ul8hiqJlpu2d
mGBut4c9QH5beojMEjPNsXcyZJoVJLAI9UyMepOLTg6j0XblmPtXVlwAfcA8cM4bl5tgsM0G3gpr
suvR4NgAVJKS5hacbu6UOPfLEXAO0/oUS2iSR6eXBt9gSufSSLIiAeOAp4EnJe0JFdp2/Lyna+hD
Qc/YmlhB0Rj+JdSII+57y6j2XtX2y2s/eSYJ4+15O3uiUdqWPTukcW2JMC3GTgEtEpZrzCDzFcl1
sOMOal13JYJ3aFPkwcqaP97Mb3mDDlWwyTvYwxQtK9xsEtivS41bMYv0Z5cS483/+zJpRHic+qzr
gC2jkGrZOAFtBPbdfmnxUHfca8Wbst4tVEs7pFkcIKLoTFNclA508JmsblB5GaWW24NkgEEalPAS
b8jEqXySsuqZGdc6FH/WA9M/Qn9ZX+JPqYOrqEC4duz3VME0N8JU4WlIaINoUso7UMQOesdz7U1E
dmbVjN+731sOnnoypDHqOxTbxFvydOPhGw0X3PO3vEkrwfarNJQSmSJNZYjFCJuFK9U3CfvvaKaz
eWI0i1gN/feax/IJEEcbKbVQn1fI2V11c4CrdmmhHJ4WoxHwnWwKg6V0ukwymHYbmE3rJ57Dff44
mkhbuQ6w/lL3mKOxJa7scHetRpJUYdE5DsHohZNM6jmiY8+gVRAIEeqC5x+nNuygiEUf0szwGOWE
TbtoUEBmWFPcoVQJfWUM5NfU/uaXRlEwNnTv9aD3BHvY897SfwWUyi8wL9jUfXpQfeCEN4ZoVp+f
UGVUWBSu/+Bj372JF/5FUBY4Ix7Me2o2lMLxraQEiNNTfRKOcvNNbt2FY1ocBFm9Kb809D82f4Oe
8u0tG2GSAY9T39SsWAkustkHoRu1BqL10/tS9qLwcq6vkDoYYqNjCD2LHXtmGc2g2FmlXaGhOelw
ieg+vB4QWEVgfUf7xmph3MR0tgsWrvMvA/iJZn//e7apd0BYzU8wJI5+ycGPrfauMIQnffoJACuN
8IFcXWRTU4rAXIhD9JeZgoZo3DWcJUsB6TgJK5RIjfgd4hYNVB2AxyM1nmXk92Uf1P+cQrRuj4CH
dII29XirOGRvfkJQI0vcjHU4foZ7i8z8TmkiY5WfAGgxj6In0OUl9xMYEB9MSqZH3iALS5ccwuln
9lM/jT7w6UrFpHwkWAnzlr903C4BbuaDkjSzV8PggNJkDCbCtsTmFQcsTFPJL9tKRSDGZQ0vQy3T
RPkyHhiMiVU/dXyuCHJs7ftjiVB3ZW8SMFCbTaVrKV4AIfTUmEKNw3ilEVCMweiBG6oOp6TKGC5q
bF7wkyqGu0CvA9nrKdlFEoMtPTvjtVo2YMCAzUcFPgswXWuxc26u1DfFrfDkk8XTSpwgh4n975oF
8AZ/vlrWHyyRhl1uR7ySsBsWDgmjanQoc8oCicfihjs98gPIfuOSAU4Mp1pi9l6FeR3PBPvwLHxS
dcu2qBRLIn62kY9QCTY7dbK440yw0d3fipW7NvJnItroOW+Pnu+edKLmxSb5v3tR1me/d0jXRvgb
7d4dK3KvTIRhIm7mjFZaFM7hO7VnQqLfOhw0mgIgC1G2OtZ3nUe5hoc6Gs7SF6/0Kc+UdBrl/TPr
JuRtpELZRma7UiMHvVnIYlw68IgXPTbcRMghm92jxs9fcnXG29SGsxNo1UwSACm3EbNmQhFfvA21
HHP+Cx0Vn421eNDHLeRsiXc/SreO6Tj7HaBTIXuiZ8XtAfRxdwi11uFiVLhb0Bnem4OstWSAg+La
FQJsOSypCDtRBPfCLHVP0RscAFYAQ/P+9Guw+/WNAVhRTmWJjWyfA8vLK3f7pMm2wOsb6jaPsDrd
X9VuYUUcBTLbiT1oYwIE2xrfio8KNzMXSj2omormi81WNahY0vQ0dW/awlYrnqiv/yHSacj0vxN9
4piird3opT0KE4oZTLpeaVFLj8ktVWEwIzMjySs6nkTZOwe/FxW0NzQ7c3z9uaVYcfQxIchYxqxz
wovK1XBnxZdzUdHHCNg9wttPqIEsHNr/h5PEcK8d7tEzVfFdMPXETBp+Lv/M2uBAuZmq+YckrFC0
kXdj7QYKAcG+eEhGBEweuLNmy+Au2qgd/mhvNVm1innawE4XKGTZ7sh/8l9QeBTlLL5XKDKR1ydT
I/sE9AZe9ijkm3SS6NQarl2XvxY0yBIqF4ZaI0Sn5ecFEk9GnU/uSEpXQDqmsqek4/UqJd+pKVOP
+Tdrhc3zgd/VI+cILZNIXEFre/ngHNzQVaEep2t70NkF+JwSggiSbLN8NTgcV1evf+b3ypAi5k6Y
uca1tMAlM4nFwbyablTxJOoVBnFWh+Pa0p2FQFKjClIdMDfJ7/7BTOd8dKS9qMIa/7dZH3pjWsLH
Ml6LxeX3GM9nn9DCFOvQIuK884LyA6mojIRqJfMq9TIo63fGXLAxEoLDthVVqAp1e4bbWFo0uUd0
NFm12DJSlI49ITbigcF5HSdqtVScTgtDGzqPwUJ1Klf1Efug/0pUSL+rTfBFHxEj2IccDh3wB+Uu
h0vc0GFUqv8ztvV4E/fbmePYfr+PkUGbPzzRb9oNTEWwD36lIKitlQVhaBI/FrhG7t8xu/hhlEwP
W3t+Yexi7Oq7OdhK5h+5dBBYCMmJsUqlWS9GoSm3hxKWXtkfjeK8ULfhf8KcbWrMHcPiHct4VQ3/
ef+Ed8TsTIuFTUJgBbhTpbmZlCZfVmbODl5H49CLsWY0Pg6ePovuDSlMCXOP/aeiqX93GAGfLNsY
pG8E1rTud8532A1MKqLZxGo6K2wueOH7THE14i7qok195cpud7hXpxHmXCJtT7uRkFOupNI3kt7I
qMR+xUGHfaWS7yCuhkvy5aNNTCtQsm/huGwX5tmnsGMtqbN0D9Rl0e6rNwJjK2EWxPjQ6gd3nY+w
wqlM01fIcQRO05Bf5XSsbipfMImmu/YrCGOHsg5HlJ47V0JGazpGbjBUldWRKCOjJanz4QmxLgnh
EwPqgC6JqDg9Nkch7A1ciVna9tqXmFgCaAFrgW98Yp6oyCJk5iSByfRde6HiMAKLS6/cd2kN4NV1
bXvvx9apR1JDKdqwWamBTQt7vkTLwW2Sk9g858ULYgreBT5l0SM9SB/sCkwx58D1QBml4N7Kyc62
ZNCRULYIwCdGc+K9KVB5YVHxD/ZC0BHcJaymMHTd6yt0S+Xom+EqVlgNG4CDFqlNlhO68o7TKuR5
rWcg4vgk1kFLjoqEo00RZah2a0X/DlEW85tyYn7kZVfRDBInorDYEsv/N7hmV4yJuH6x2J+2YNq3
xshq8YHVV70Yp6aRA4nClaa2ICcSqdQSNayjNucupt1WFXA9CZ2uBtLqYqH7lFmmf6AE8p8UA9i8
Kg16fhksM7dAis2CEOCrrvB4b6Ry6ZMrq/nYIkIIgJ98+0TuZZw07CRaPI04GNUlWayxHFZRcSUw
cQlx91ajB6vSdKr/nWx3EP3JNkYl2RBG7wJy5G7ssh3z+WwRL3P9Chx59YJDAvh8m14sm23ezbTc
Pezts1ycYoqJH7G7jGS+z2S/SDVorGnPSxcpsSqN6TNuzSqwm4gEGD3glSLjLqRFMRdYx9SlBYCq
Iqqdac3N82ZoRnC1NdK33t3HMVEY6sKAjJK2Hh/t9mcI72gbP+ZjLpFbcb2gp0eqr69Sr9jLkuoD
3oPnSiVDkA0FqeOGb5m2qkq1/4sn2vj1F4Kn2XvKN2mL8cQvasvRkDoazIoD3OUic2TGg9XMurtk
Q2OsRTllUY7QJK5efDp9+Mj3oyccZQQ7h1X8oMjI1znrOAnyi2ox0iOU9R7PKWyjg1CpsDklTQz1
77XL785rB4jInjzGyllelmHgYtLvj2CxQgrxdQPfIjsEwaFnaAQkaJ1Lp2V/yZXQQxyXux9CgmVZ
xYUXWXFXgqASV8RgwfCeSPgyn+yY874/1TIgFAVZvXG93G8uhp82Af84ZKl6HL+FqGRnJFKoxQFD
j7WR/pkcurz73t+zO3L+8aM05ofjsLSwe0H6YothGM4a2kL90FZQxQbFKUx3FuCSr05yPlN4O/f9
w1XMDJ6M81pQzs0V8ixpgp2UbTee5LUwdrP6DAjNzuVQg4G7hUDYP8GuepxUUxe0Ijolyw6/aViP
EwUcQ/lrbpHnlAnV4jaG/pBAfjK0AYISswv/YqqjbaY1kdA6FifllmHaGXFfMGOZrbb7Tbvlb3io
KeiVcnGPdcF5WL+gpYOaXnu9287fZHhe9/Nxg1vqzgn3JQopcvgQ/C8tpkcuQ5pJ3sqJfA6fAldr
bM/CJFlrtyCXwLEs+IhLH9O0EABMrzRngvWwJrGtuZ1eJm/96S40MKJZQBdHOyhqkXJEvEJf+CD/
znmlZQOXncuZNALQwYjsu7S6PWau6AZ9VYOP/NUbLta05KcfMjP26K3imfazkqliil0UHoPjqKXY
IyA2CPmwHNKpp43VPH+2ffAhQSZSEONggzYOEhGqgeTkcf76tRCfiFdE4oRv8g+bPB4XCHPQPbK/
jHGgteaiWt0ZK6+PBUSeNGwoULj703S62Fv9kT0g4cMSDbfPixmmjkVpjrSE1k03DDVFJnMzuSjO
0VynZsVd9jIuJPZMNav6dM1gL+3dvmdj7WCa7ogbEoebVjqZWcQwdl62MjHSuiPCc3mtEX9yS4KL
sAGxwTlVZcKOgNz9BYzzkufKZ9BiwGtvVO5Ckx5KMDqz8JjXz6PP1IUZE/9X7TaaTrzSeeWL77ml
kLc1eL73QgtemDkvhrdCsVql7UzAvQndV8MgcyCUD1NcdN4amQmH13W6bOv8x4gi9qBBC1FDf6tb
XXSEwzh5a7gUfqHtIm39s2miOqalbvwYHZdIPJBcW6h5lvZVZsdmOK5Fie/hxtTLFQAEjfX6PBu2
sYOU/j6KZYeZdrlA3bm7xnHmZJ/6XqBRnHlVdR8QW1cKh0yAvPCyjJDuboCT8tQlHb6VlfKt2ulG
VRSZ+jn2LeJF2bia7t9ZElelZNu2PYPkki3s/CQpeMgneZ4480BLtOo/MNt1LXKDvvd98xiGoXmq
Osar5RsKIjeTbnytsQFCHEL5AQIP/VSMgr8Te0GIVtB9C5JYXaOs5pIW+ZAdKfCrJ6RpNWA8iqQq
N8pgB1CVF2aJr1QEZe08MHX3w6EkkQtbxKWtEQcm63PLWaYtIDpVAaQxmCT/yijEyjuipVrO3//i
jGVwQLSoZWe6q5BFx34wD1vYSJkkpsOFN9thm8OXp/8N+YRzcPHK6Euj6pVYe8F/DOEHHmq1DZ2s
8x9v/OnqYRbjKmrdxh1HD5ELTJsLV4RyIzpslgMJcSgBT/cyFa0PsqbiuMT7UAEh2lK4I537N9px
410OChTzm70oGtvgHQxPjOoBFlr33UVqzGKI+gHzmEZdp0uWdOt++8X2UTBLAY7zOjBKF7gSM/Uo
9OuNO6pIiI1+LCg7UvbspmVJzXthaKkZhumM5+n3iDwMecGOS5EnScSVCAZNPLoE9BoxV56BNGnL
rk8R1rdA93nWRNM4CJHKsMvW87GbLq0ZTJuK8slu0SG7eottzfhmBrM8gXHf7k244mr7nc5qwG2B
GiqFJkGu+Br+NcxGEBlu4PS6onP+qmRwd2lq2QQlJgExKLrvLQG06lY0WawOWVYJ+h+rg+/onjCg
lmxdGbUC4SU5DQC6P0SDB8I/1MbOVrpDniyfXoUaWN08uL3mZPY+RZwn2d7MBnlQ7ZnA2+CUKJZw
6b+YM4+xvgM+M7c0Oe9cYI9ieyMKnO1pAE2Cn0y7+cnwJlkPNFnF48MOD/LWd0F7Q7jZG+fi3fjs
ntYKTql7twRIFfSDYUREaATieNUkNy0yNs0CPTpp07WJCz4u0A60n0eafq+XJyrtiXjr8j21BHzs
nWfmBBTz9AVTBUC5Pu5IZboXsOkaSVuOTRmFMuA6i63NIaN0/WZvXS2FEIgNHB++txv3QG5ofmAI
pDheIYHe21vqVnLTuKAXGQ9qwdqiguWXINAt26onqLEd3QGx2prcr/48rxwsDroqTs6hSK7CSmBP
Xe9EWlg7ptf/Oh4AkhHpW5mkHj8xqXXgTsB23O0maanSLexGs6YMTSPnSzfaUQ7H5lqYsMbCLPAe
NQfttB4uo/KCSwQaceYStB+r0QBWKKn7UhOpAB86r5edTgvwLn1dtdyWEquQ7Ff8pxyrWJANc+Qu
WBKR7r5SEMZ0sUewrF+AZ8HldJF/75v9Plud9v4QXMuZ0Sec8WCLARpy0psUDdT+dEMPio6SxKAY
1VhOffuvjDYUL5B19AVfCV/QxwcdPzBp1PSXkVmsmIDHE/1vBJv/YvyYUSGfi56A1uJH9Y5bBLow
uigXuqynVKhEMfQJqmk8Y55H25epGIuF4ECevqe+aMzCFzZLFORoSkGmV2nR/AFgTDd/YHmAGPMc
O/dFte5arOLIs+NoXJHFYFnI1m9+4bF1RlwfqtGJg9iiot4KTFjcoKiPGFwMbz43cHkCrXYsbs6v
up6dO7MZHt16slWqdywD5848m6sVEDX82EJVM6arn3Nu3zGRM5obY2T8bxbR6uznZuRo9/EY6fKN
FpPBf72TRrXG+VuAWLKVECA0x9GfckfMcdY8nBzAxMoIZBkHnCs4c+dP+uCPyaL5zh70GTnJYqA8
VNUdc710WTJIb4EEngvDcbj8fCJfwHXYM4UFa0roZL9LToQfeTUBv3q6rbDR1NbjjFa0qAF3mxoe
Uz01auAa7CrLCYaSY9h9Jo9p/dbLJGq6H+zcV1pfwhlSkoQaOkpArGYJ+UkmzJVoSdtHJ9BEfzTM
LNYUR+WqRVno8DOmXOtGPNFmhpsQ0mRskuXjwv18vUQWSV76guONsOhSROdhlUlGymNX2JiEvIc5
gsECXKLMF3bNAQA5OE9ld/lyWShqtSorhUgXsp5d0aGnDToByi1RsCrVPf/lQbxsxPCRqf78pm6g
cJAq+xBQdyxeJrUAJnnJ4brLrVqlWmVqK1sk0xqQZFRFSvoz9vj73E2XchMvbOkdw8qSSL5oXSuW
7z37HxvuYNrX+xQNED/TI57iy3MBoHW/4h3KSawVMhp3rSqjT2f3dMY3qBNm5LIgwcqXagH9ScQm
J4rVBvGAj5ojnHYOJRceQrKH3aYvOpogrO6fRz+QeF4sAzaFAMpXBS4i9MZddQyDv3s3ituoBggs
twLl4V8aHshs4MGqgtUQYA9Q4ug+eXGK0C6C5q9cobQIUiZSHektnFv8vCc3/ig+gtlBrr/YsiUk
nmII0jAhEzrUjb9tvUJaksHiR0xWLmiztleg1KOjpA/1FSUgdUM9jDie4Lo8vhBmH459up2DfKbL
NPYsK6qT27os763OHiD/cFSAjiXNf3UzMA5bxDWcWirlhQcG/ngdbGCaim4GW8JJRzRNX2jrwjUB
9CayKw7GDrOnApu2Nju7bRKq6ftfAObilnSPcp3BvnT1tQsc2CKx5Af9W+xw7/k6VzGKYjvNXOYm
L+mhV4w6xSjtmDi/TWFC2pY3whhSTqeuWgGVp9T0KF6XOsmAX5vhXPIK7G2/OyrCoDjGMSKXi8Dm
puzky2HUoBhPKWpU9X53y7afRn+2RsgRGjJhQ76FjhLYPSc09jrfKHIiuiojeqpSA04R7gIYWwDP
5cL674fnzX96iZvhz3mP1hDj//TAZRl1itfkABJ1xl0e5l1ftihCAiB4Ov9NQivx10nnb+k4UJKf
fz+1ymRgPMwSEjHjEQnxX1bOqLPB+ec5YIoCQokLHe0dNzmAw0VomLNRFFSjIgACZZfE+NtUN00A
7l8+4cbkeWisb+fk8t4OZE6g4snS45sT6yErib/soc9oeWkRRuGsCQcFQVy9OKa1EHZsqFW+kwlZ
Caj7X4R9YlQCnKj0uJhJlN5wXKgRmlMu7yCxUfBX89V9GKLavfxaGhGLvpMPmnBY5CN/A5xE/45+
6WmlHr2qq+zbnsu3Wa6vYiaJnm0Bqh0AgRMEklrcdbEXKTd8auiqpt3FWXXTkeENFCca2e1Rkxvr
vNYD2GhsDb6ymFDwhUnfMsRyJikDuF8kl0u4YTDOKQ/QSsP5wj+WjYYnECJ2t+gb9aPHE/PD4f3R
Zl7k18uB2wbTmCHrMjImw4lgTlioGWxW6kOg/h3e/VakqfZdYvXl2HDRrDpb+BAsGmrezyDnZ4hj
u//RGQer6exB0vtpevZneLpve022PxPbwQitnfX5NfCLaSZQJGWTJ9Lr2nK54IQJJHzdubdqEvLk
BZmrR91aWCLIKnKKExVonFhFWmikF7ZQ9Wao0pRA7VTUM9NT/vXRU+TOXBeyXtgeXFjaHwoQ1s5Y
AAcp8rM6kCTuZx7tTZ+LCHhHnr9moLifVWreyNphrNvQrTjw6ggK8WqPGxzMYG2crSEvUU7f2f5b
wZIJF1opYKSBkHJqQhvyqAysG0Yz7e7boEFXLBZ1kSOX0W2CG2VkphR6vaQouhqYt7+/GRokVc8G
gO/BXtcNjeYVB9z8L+3LxRVEy4fuDjyOthlAQaC2DrNLJvaCfaIwqQs+dugEVbRJYR7reRuJCXB7
OcaPVKYyQwG+bD1OBRXQWpIhkRr/UgtpDT4fHnA8JOBXZ4PYSLIqFUI/3G09pEuC5cvchZNHXgG1
+4u0T9BVq0YRU1JPK/fUREos1UlE9m+H73gsFn/iy8ZF8GH7ZXGUai1KvTlY0skWczJpE3mfgLzR
+8ZWGXNRmMG2vpbvwKnPq0ei9S3hy1xdcMyD7H0EPsEu/P26Ju5T0/QjmVLrAzyNWOUJB+RUlOjb
Ul/EY6jQ3+3ojyM1PZeXOkcoKAzn1bi26UqIy8sNsGY/b+ddul+3MK7Q51VFNxNiydRUxKiqQOir
oZDLD0poq/lfDTqHXMI9P72nxNgVVmYAJB4kE1KJ049yZ+CxybvShQ0CvazICC1D6aJFxLZFzs02
McjQeanZ2sdeZNJ2fNln4uLbf4sKcmFDmLww1RJe0fITFhtJyQzmLDmkPwLBx0zv6ydYVbO03xS+
Hp9W6QQLd8Ve2c/0Hb7/yFGujsreEPuZyiZJDhAM9wy3WAPWfYic3N8P9Xal3zZW41IaQ37v+GqI
QPGn/6WB/nsZ9SegCnfZ79LYfR9hdg3swqb9jfPTM7RUtrYIK4uo2pasgR98+UIlmdHIZ56HZcJm
GVxeqEDwQW7P4OSIqxBpAiVE9HGY+esreVMhWlEHGMVXw1dnPiYmC+H1OD5pa4Hw+cg6xM8/eNj0
q2tFeyYHKjKeGrWrv5CSmlU8cTBM96OEGEge2KjQgvirWdg+EBBSK/FfM417uSyBoMy7F8F+jTHB
Uy/9nr7EjK/Q4raV/hvhW8GA/Q7k840tILgGQIzqvHPjaH3bF5bG40fOlRsfUubeYPxXjsShoA4H
vPoDR0mAgNPh4zG7S2qa1o45bi0Sr1ooCsjuKeCMA/MD4jqryGEuUJvrwoBSMDGsw69pz7Cy+oMU
2yQCTblS0n4XCbl2cQS8a7chsmCu0GiRh8D5QpBzVMdbUtzvvdbZPSmP51d4qDlIKYVPLsWPbnY6
mjYyyrM8uoNwNeKCPtsB1d2FNdINkgoGkX/5Iz8rwqG7fnjcyHjrtzYwfBQpILQqtZhBWrDT1OSd
xYQKE5OcOYUQ8WVta3GjtCY9J8lmzS3acNmKuujUtC0uSrmPlPKnCbWC7eIELh3iFI0UTp+AoAul
j1kGt+xLDOsg3xXqWOmNjqmlj28ZVEu5rUS18XaUG5ZAGRCY+68ZBQOcZZ7lTPLPBe2wuDkc1r6y
7aDjAVu+DYxvLGEoIyFj0wxr2MdU2vBMN0inKGSSeptkYs4aqbm8V3No8bbEa7SlYyp17Y9rkB+t
9xUUzuBWqarlxOIRfkfYmq+1FJPRlFtbusDpw5e2QS4G0e2mAnfdn+pa/vTlVb2GUqroBDEisr+m
sPU2H5C0aaOf48Cd7NrJprEFG+QoLgIEewLH+MHNQr5PnVIzjy1cgrj9J4XTwDi30g7qiNSUsk5K
B7GLta5bcZTNGbemcnIcQNMBhti1O5ajqd/0igcqy0VmGgOZPDeAX09ZQcCbWTAi0jSGnhkIsT3N
I0y35ZWjInmolAYjrJv9aoAXGC9Q6Sparpu2doUum4V8NM9Nfx4lrk8AxRwQpBnbD33OB8gCFVVr
r7TbY7bLjDAthYo403fR0ZA8p0j2Ig3wHVJmKM6XdlkgxE4u49ODSUFWE+7M+7bYEKRQol0zNbfz
6IlqVtwkqcndB1MfnQm1O22yqYmmJdc2eFjjzq6STjYTUNyy3TRpBLqaviklw5n5FzXKivw68GwA
GKbwcInMQavJECYvbjy6cG7OLpSA82YiUhwGBlt3wNth53niNjZDZ67Br2FSIhKmKQfdSnp/uDVB
0p1yCMq8G5e5y5VH7hSDC6vEb70wBPO0vAbsxHg+de34V8UMyymYHzwmj0vsIB8xYyx3F3moUFl8
yCWs6Am7DNCZ7/vo69dUIqoIsOO0BjYeVKAxjylaupdKAf/nQ0U0QH7LeiH7jfhM5LgRxX039kTS
GMHsuOoZ7y2L3EHKrXj5/Kq9ReyUGXmvzYzhl2EH1BR+TF8JJOatPgHvY7LMuCGH/Ame3gYlE5oO
QdGT4MSN/PJK1HA3luNNqyooIx5Q/zsZKyAU0iWzHdXAQwXOm77fH8ifZLs3ghSj2g9j7rorCinh
OFKXkNlNBOBAZvckzzrzT/fjnIP6t59QPnmoKn5Dn3Vk1A5psOxSIdGi0/FFRkmAJoYPFcBYk3yZ
d6JOcR+TkgwpRwsqv7BTfysVA8lbCyJ1dgzCudFof0IUpHi0WUoP/Ao0TXxJLgT16btlkCQkyFML
mf3h0WE6UHq9rFy7Bt2QF1OZYQKEKPp687USHBDyktL3HET/kjtr3NlYaHzAjo2JRoBTgNwp7Y9s
0WeoyBIlXIG4OLT4VOfGlrL70A/VuczmCq99H6zdSTgDF3S0hkAXDNDqTzitK7bv+x5tFyXau/ZG
Dgv1z7Jo8Y/h/esjP4NMYXLTLCm7zA+Hh8HgRZYD8PuRktNmt89U0zjx22azRVHJM14p+kE4rep8
O8Km1OsVysanmxAw0j2baEkbe11YOmju+b/bDsiiPUuWmMw+3S7XiS6VS8m8m2ngd8mns8Gt4y2C
Tk73mM1NHuPmNSI/8EEV3OC218uzWlXZleWP6ro8ygNXJoHLTMS7wjwGGYqWH0U7t6nKBBFp41cf
tUVIAngGTs8WYVPOzKAolDnru8s5bk8/EoXwsjh37iKACt1I2CN7cvdo/ZizHu8l91jGfZjHikyB
fpQoLHi1m4p8sdrrY96syKgiemIrT38nZxMZKVgmxDUFZdu3zkOl/9u8dNKm8brnBACK+jlqkA4J
YhePGOrxnGLfzDKwFYSQgYkkOhCnX+DBdHkWd4VZ/f/4IL4sD64kTgIakeiRU9hvxKM+ssXfwC/K
8u98bLPnky23N2zLebf5CGBYmIDHE0hIQY2VnA1omgiqI07UdUfMJn6B9lhVCEG2VO1gZYFcUDFH
KF+3nTYpKMwUdIJK/loMmPygs2GkzB6QFDvJrrdS1KmYfnBdXIjZQjxjiuRBIRopKCcVXaNMMohv
LbObYocbsMcQ4qeV/IW8qsQS4btcXOguZ8n60zVafIhQbGRKmBPR0onnCVt5h8ncveHC9P0uqnjX
2F1gt5wu8M9MrcpwIjV1Ff6WCyHdWjP/TSNSJoZWZDKt+vNUkK4MHBIiZla7WZ7+DGWwYRGs6ulG
rIYbmQng7odCZC/bAAEEaPO5xLS39nA2tKAQsw/Ahgu7GFfnhVNd2NENSjedCjTcnKiJzadkUtW6
t+l1N956F/8Iix6Gps543b5QrrLoXd+aBQS7QqnnL+nB6MzWLXmzLNcXolTP1/UpRUcYnxAFotMw
MuXX+X8BX6SgRN0AanWQXBgVbnLdBWwk9SF8KzBe0OsHTMgZq+Z98cbphpijsVmDK8//QcZH5B/q
TOP2Wi7kSPCUYJdn9HOZ0Nkh8gG1mLDR1wkHLg9+FnQ3BWttzbE7HNUBgFUGmo3zHFu1r9JRaeEg
q6h3hQ6clb9owisvlR7enzS87+dwE3UxJwRRePQVhSx61DOAC9WY5BuaIHaIhORsgcRcccECVZzr
FjlQiJpy8uFQnGo+09P+WV4MKeJ/Ow985pbc62EsvIGYyeuZJNbvKq3G4hw7A0xrPePa6XDzgLGV
pxPk7gw0zahlJuVx1Z/x32ylPEznATUjja6GI9Mg0965eWZZYQP8dxoY8/4QWp1dUR+5Z3R7p2kv
Hsh5gVJt5yFx/uDC1cep1vVMvorue3Cg5J6d74sl3AovcGtsiKRWU0e9kcEJnlK4STxiAYDtHB/E
wH4LMnndCA7UGSu3NvIE/jxnD+mPM5rZ2IzU0DuAf0E1t0Df6NY6HiwqAERP0h6bebKCNRte1oWh
0+58PZkrA/Uy+f2DxTv5DGcnZMp7xhVuIJ6fIY+z9koCK1PoBZhS130KgYzMNE+N+QOmWp5kjwLH
lnfOJ9uAPjQ5zsbUhsg1QwXFYbpBl/1aPAZD3Ra8FAxlMnVMxk33iQtzXrdFPemudiJ6/Pms6AkJ
Fq4Snl5DZJerNOH3ctum2ZAqGQZa5qxn8frckoIkOfswaWxIWS96QvQV5hozDdQ0Gh1/i1bulGiy
97YuERJvgRmPdZGab1WbeRPsmEx3hpCzaQwbAuwc+HceSTUKHNpOgFxSi1JGZvLBKXbovKkUMzY/
F2lRIfXzOIPdnB6Hryrx97BA7TQeneJ35mxClS2ww6mQItYWf3mIy1ukwMBVxDCAA0DTbthkhjsv
O0CzAUMRUShfmSnAYFWmc1ur2TIgnOcGaz1B3NvVrw56xiTO/stunXWQ0peBt4PdBhOcSeGj4lGa
am1H3A3ABF8mXcwDh8hcbC6WYfVIU3OUvp38kAbjnQHHHYqdIsG5UTra63bJCDyrSjozI5Q4OBsC
XUt/1HcqwjgTyhZd81lpRu0wdUPP+Rqem/6407elt9ZXAsM3ZQ17T8pwcdgahlJ8LKWwXNvvwVXR
LEyyRpCfM6IDkOtPnTUADgpgVMUH5/St2A+9+dKCI2cnD1fJB1Cqy6+UldZ5L9AhM9D54bk08NVI
qGvkW9/GyBqeHvzFc/uXy+a+dNrTrvt39mKZZv/IHOp9tYbiHq5ghgrMetqy3izqcmDjbB8XWXvH
znSPiapD2MZWiSiGLBwvs2/T6dm/FT7t+h0ZJi5hYHkv5m3+Maz4fonhDthiqAZ6lx34sNRKr1Jl
TQOgMhNvtYJzDwzPBe8XFc5YA0nQkCb2rQ7/6f3mJ9uME7eggTPAwxGgmUvQ1sSLPaYAmjP4Z7/u
+feXtCnCZQosBS323tBCPyfKhaxJsHMyqUvBU7En1iiGwmXNQjHQTNkcYsRYc5324E0jvMbXfMWn
cRM/58VsMAJPWUH55GeNXPws9sszhvbuwdecoJHXQ3C8D0aYeDGI3BxvRCRnu8LBw08RdFmFATH3
zCFpwhsvIJFDmfmTdcd0KTKGW/UBKGj1r2j2oHYdYtJk4z0VVBfO9FPUxaUj8ksjPHmMBC/c4a//
Ke+GuvgGOt1LciayfUPotmzdm4wA5BCzs1nOesVPAJ3wwUXBVrL3b7rjn2ha/4uVrHv4mZgIBWep
o+GJPhAYLz36/WYLjq0BqjxFtw4iZBCD1hsNUaSvsrUtNV8MHeCYoypvEKfIip1UOlRMIcf+iM3s
j6laD4tEu9Zy7NXEtGzJxv4VfxIcHqvBBB3Uuy1stWUGsi8kSkTmCtd+Rs4Ce/HwMgn+yhXQoQQF
tpNw9u0BwlUl9XTPrybvrgJ6Pp0AJTmkA9jj4Kj5QM1DwZoUHljNMQR44W+PiWCx1SeQyPsA4phG
sk/PimpjCBZvqQXp+CPIAkMe2PEQewK/Np8XVinnOSN9QgCfejXNHzqo+fOGK/eho0ICR30YLID5
h7E27VttjSK2VniRbOESZrqMRqBM7vzCzOM/DsXaGOhIMIioXUPYlkOYg3hGTTTp00hvFDZeUVL+
1cxgpdkZCYeWTpOBLKkiUIzkm5a7iSAUQpIqfqcGO7RfoiCyxGE3rBIkeR4wN8RUhBiw0NEkJkut
JrGFn2QQyRHBu3o/wZAX2fwdufSW6DYZoB6KustzOFzpQMS9RbcfzPnueesH8a3QGMS8D/6Mepc+
EEoL7/oz6z3D3lggwsvxu7Dg+eLv1rTpbdLA66CP3l9Xl68DfwTBHva16V4xvtIYyqz8PNeJWY1I
9FWWdcgdnmcwuvJX1ljUcgMjkGUoo7iK2bQJtn7w1PfM5ArgbFCD7CL3FgoMaJG0lRGkME6YUZ3C
KkNhr/6M7bIG7DBz3LzlotNgT+we7ulmTnGkIRYHrm7FASlSgNXhK/dLfWdJkcfVZxEDmM5GVi9o
7IeuuyshQAGDNcVyCRqgZ0qGO4RU8m71h4zH1cq4oxddp+hELhe+ueWetTB3PbuL+E5oa9WzQwZq
FFGxtunt/IiqdSbVjzcQyU4goSjfihr0pynpwCQ5irZyIblVOvTuKDnwQMrXVyseUKpt1aS+385O
9qk+ry1+lkF5fqOFee/Izshos+y4kiTcUlywSj1uVrcJdL4vpEvo9rZbtddJjL+b+TProkaTHUqv
8pMEzIQN0RH5bL31dcewojyaQdjoSbuAJF+V4iP1SMBMHD1U+NRfsUVDXjXach2jcT5P9kh2PrVL
pAxDCY4wBepK6uYn1XHkeUdDAnJiSeJQIAB1TUbf89xj1JVy9jS5Zz0Y3eT3vbl+rjv+o8N8orzU
e4u1t5TG8IAp7P7hQ0fJgE2iGUDV3DzsG/VRya1WAzWCLqscmGeNaXvFnpMg0/F7mD5DN1KhEyMP
4wApCZ3wtqPiDU0w+1vHRdCGO4IdNALnsuGg9Em8Hfd5Aj4cmTjGqLVtvLFOxRtWRk8gA4h22NJm
9FYurEYesp7Z1p+79FAwHl5rPJL069HiKgEikB+zf56f6Q1PB6x0zgrR+z7HQ5ldnSfX1PfXyrOQ
pTTknRRPkoIdbak8yGtbeGL1yva41wVteSuaiknmaFy6JQ0tBZLVk84RX4Mi5dSHVUshsBTrWLPe
xxjdyXG8XSgZb41Y068iBlfBfodnEhfLQbsr7paI/wKrRibq8EUU3FyLwSURwpz5kIFTqidN0x2p
rzah3KEht2Hf2EZtkyNI9fMiluYg0dbx89HxMH0NIcmAODfFwQPUt0SfpyPvSeqHbUXibBJ4QmW+
Po2a37lawXDg/sp2NfGxEGsQoGNDljiwON3y7p0sR2sbe06e/xIb9usu8PeXXI3BO9jp/f0jNJuW
0IbR8NwOYbo4DgZTB8SkgCw26vMqNNvyiEaS+XFpTLWFoVmlr0f/mqScOOorOyPo3bsIKVdxSae2
RWWcjxSakA0Q0+7c96p9aQjEoZzqSwrDyr5DtaAYV25b51/74pJGeIt2qaLGav4DlDCVRRDS4Wes
GHF4EaMzGYVVj0lezSxTx4D2S+2Yd7SJXL4A5mr+U1WPwcTlSDnD8ljSQd7C2w+33ufLXcjjxw5g
r/IboA6oiIxGB48wjKI0xkKq9zyysyVnyEt4AxrvnUO+8zb632otGwUL0SX5pr7dtv5Wi8fWOzum
iW/UPcwdllkscKjsHVH1lMZ8mP24NKkXW8JHE44UF03f+V+1BM0arLztqxJ69j7atwJzJL0KxgQo
2b8rNj7g5fPZtG855+/NcvyX08PwKjlFVrSkWR9HGzU8MN1WsKM4I+VVYY1g9bQye2ZOmLUg41FP
CM5Jx7m9fqp1Jx95nxuW+c4pUBA/OYYeNfr7/wAbZYhqfegqo4+IBs/g/UNmTozT+7nQ3DQYvEkr
5QTDNRku7H+4H5Q+DJQ/7K6AU3zxqwYx1ONE45d7zenJ4+GiqS02W416yTsN13GsdQyX6BOkn3jZ
/zqwu0ZQE8YiG6pGwOJtvFdh7zlyZmOExHMd2XQ7y/3UYzwEgBgYm22yGSR7u3UHrhjLIunCHvPh
eSCNKgP9aLzjwmkXQ+Gl0/bgSZV/VCT/56cELYp8lji15guSOEYUWg3Kg8VvBCgoswFn+19Uc1S8
/GgtnRjcbBSfYD/Jh4xHsbRHbSAaRao+0B7YvalAeCsXOx+RZcJBTqgpS9K8ps/nsr2/SsiRPZmt
WzjqQlybHSA4GjtHvxOO7P84VUBigVpEnp9hZGYIP+YypZgsHcoGoh1iqDCYQGLShqQDGMXxVN1V
1DAw764gcxKNyOSxuDjV7CkqxNSeNMgo0VPLmW1lw3Ciejy08RGod0EYeAm/GD+zv32hjSFLlTp6
uyjGVieditmysxOITDq1xOfbvIfK6TvbORo68+Jo/nAOCn4bBdP3+e4fz6s/G0Ljqsj7GM7SWY0Y
LkqO2N17f30G4x1TeB1hWLba+lxu5pOcGbNmvTdAKJC1I22N4FYy81abKWJbubftrR7JxsGRlOfh
fl16oQwWU0OkGPVW7T/njbJLSFLJk5aFMvt24Nd7GkgIWV9GidGUKe90oVOqDdEtPKRH/6IEi6Ce
8ioOBvVJQJbjRBctSWYVMIDHx3tnVmtK+UIZBlGCZwDJkxC4WoPpdsbX/i2IH93bb6/W5HrJ4Ukd
nf2/TlbAxf4NYjERYNShvhlg7Zbc4LO8/Wy+p5bKgVLYMMr31HKxML4gHB0MKXv5I7Oi7lsvS3jj
G3ybzujtFl45G6Lq8LFgzS1LajpKZ7QqX98jB0S+bHyVvZsFRGeS42zPJBWkP7kB28Vf5tRF1Kz/
5GpY5/z54U7TFGIZgrwkzdyZCJd6mjq0NKOys2AyFqoi8IM1qB2ISWkca3IrTIQSWTS2Z0jOAUdU
ySPEAeGG81LMFk48XomBfM/iuG8mkWVTtBoRaaikCzHcUUzOjGPdZBaw9EmPei/CO0jqIqfmoECs
oKLFsYo2eRc0W91LZs6iCVQ1lDX0HcP/Iw7/CHa7H+kMLnRnwtjM5G4aOdbVSnVhWFWxM4YW5/pu
EsG0pPu5zZue69g1HsnWWOd74WrmsNdWyGcyeDN69cUhNgPhVXVWfhiBssPOBcomPSq2rkJDVwrJ
SxYkb4Klllx1Hl6uzrFNivkDo1i/qVP8nArcr5kYQYht7xgdYowsm/WNevAnLNWW7Yl3ptc5LijL
/5+11Pujh09fCxZa0Z9EONHptKO4xQOaNM/StRLwAQo2f/y0tblHhX2Z1N3uBF2RaZNOXXXd50qb
kfqEKo119ND+0yV2OszHAu8pihVuupqpvewkxemR6BKnhOQcDTBWKzxMgWtFd1RrAjbhPCPOlTVS
+L341bMXzX4onmA2yR/UBBe0TnZjqo+cWNLKwCKE90D+ldc7kv3k27X+BpNSVGMhlOy1ACrn2RiJ
9Kq2zPB9dwpNvKM5S3zkbgGNiT4K06QmtQgYCVG3VxGOddWYEW86hMnjqWE8wlyqyMVE0V1jV0lM
05R+mM5nXo2aXnrvxRYgpueZbXA9h/XF91nOryqwElhWh437+7dql8lfhlwUSqRa2CsmLq1QWc9A
egZWCVHAV9Bqn0lDVt8NxU7v4nRUwO8RrPBLqd/RZ4W0DS8mUwLun3SdFKIzQeNGcy0RlphTUoN9
GLnyI63LYfXbBFN5ywIHztOFwH1rteEE/UREVSHrWQ2O03Oicv/MLw/Vl0D/86K1GQFJipHpuZBb
UomxnTVCzY09Qf6m+V9644QcpWprdSCzaHGEBBrc5Jv5lbq/JMsoeTedM4gaWkf+0TncnAPdrlfp
qWu3bSWoH9UKMw9qVm5aObaFUXnTyNKDZPaaPjRx+HjTag/bIefpwYqShklr9pGv5kEp7xmH7LH+
TNxUpy9g3KQropfaQ/bxvLV793j9B1gVU6xchTrbC3QIcUTM44qSNkPPCgZPNmCeQCvRxufLRBtx
/zZv2XSYIz926LNpKsrW2HStktRVPEK45cWkUwhaGMTTZnieVB6Ch3yNqr/ysPMDatdb/FUFpbOt
q1fhuscl2TdyoM4yMgPwKrIIJ1faE/6/NUqJp25GYR6yhMKWmz08+XfYEbUADCiz5+cZNCjh0qFo
ZqqSAZzzRzX3aBhoXCsBGsFYhMm071A9cYv8vAApMfJvxMdGi5BdbrxYv4Be1BXsSmKRKE/yrrrM
jVNJDwzTF22ez23ghcSQHReEBHedyu0TvQ7rBNri9gysimS2h7xDHJjIRZz9QrhlyXkCcxm7d0W5
Wl+xa8W6F3MP8yy/hrHMf256KLCNt8mo01sAC9eVJzAnxN2nqeLg6tFa9YuFRgPBPeuj4LuM3VAs
3jFkiNd5uC4cxbv/V8dFvMoH6WddA3pTBI8TcGPWFOlniPdzBz6viWQuxU6RYsLkB8nTqARSiwHx
B4Z9I6FmpbDLNF2X0rUjn8BBiVSjTDThJo97d+Vn36FDSmERx4fGyjGH3tmi5n5mX6wbOpU8Ms/F
VdJGljmuFnGhpokBR2z6bweBvNcQdWgnJHjKVEz6ynYSnwOVQQxjBswyFNcLsvrOc4SD00av+eMA
9g8GKtt8IVqIRn/Z2ZCEUVxpGzrOyA9F0F0XY9pFNiRgu67KxU70kwa2eqwRO6Tv/2A4HE5GHVDP
7bluT9AEnKyMsDaieKWhtY8RSkh+ZwqDhXZlddJsEwhtL9eWsmG8HhTg0aiwfMetGDfQTyysA5EC
I1wxXY4woCqqtYwnN5EX6z7I6u7skmrQ51xWYsbVav/AWm1HrLi7WNaydn5r+MWv+KBaUYTO59f/
iilGfTRwlVkw15XZcXpvOyTNhs9wPXqKBWn+F35X12dZgEStZgDvLhNfjAFLmFd5QIA1VEDBgRTI
dzdemhxU1e9fvq6VXrFLaXJuHAOVTnRTNVImG8WPjmxLtAwhI0RsWj0N6gsujZFzbCG8nMp6J+ZW
y6qfEikUEtqsWpCUIadEzCmRo7dijNgC5UO1NM5+pYbJkqRXmp+ZJJv6uDhnnzPi5GI0ZCajgAp0
067cm51WHhCD8ar7PeM6+n7kpL4p4Lp1/vK2ccN92mKmZSxCKxGIsjV9tl7NkfJNOBJYUBJCPs1G
qhxLjVOiZlGHDMqcGVoEqVmz2X2C/tt6BLjTypr+rnPrhb6YYWXjy2y4pK2PVq+RFeyGAVKfm2k5
gCMCDVDvLhIy7DNLGRMUVCFZQInduTS8zS7b3u5TTxYLSakoiVxWVGzpD/jZAfrS0y35sDkyogLX
gMpYzsd5TNsvlEB88ij53eBMjY9aBqDfKH5XNSSeAVaBcjDmhuT89IkI/JQwn0eWcggX0OzFZbW2
y0pvStpINDB4miozvngyECz2jq7zq1IbehIwoaWas5YpqR7jPxkiCNrI0b7467leGfUrYAU8V1UC
LWy3RXkViqYYVV9Dn/7SknbMvv/Q3tEzX0FgaLEVlxJIn+T3sqwNJEA7AuA5eplFk9e/QGNamY72
oScezNAfcQcC2iJVyHWEzRL99+fGF0XcmM6mMRgQDYfPcdAP/mgEQPTYRwjiN7oKtYAlCk5BQl7c
aHmFd6/rLP7WmuF1NEBx/3X1gpuh8q8nNJOXZ6uI2tOw9qqkLIjsHp7t4q/iW4+ygzRWqTq0s7HN
YJ71GeWeizNV/cROWGvilMDqP3haDc/CKWBp1RB8G8hAUyqwcQuEmRziUKAhRmwIB7/2T14K7sam
KCIUlh0VPg+tVMEA+MgtyGzWIewxMHMz4NKCDtduwwx+2lG/XJgptS14GjY6oIV84BDHb+M0hss5
RE+1in9r8auevfIxIPaQJ2wpQ0ZwGE/a3KumfYeN0pkUpqOml/T7fx9+s9C5pfy3XZT83kVni6EQ
Q3+EpsdpH6fyaYb8vSxkP5wKGZ5qVuFaeT7ZlW7OF4lULA93iIoSB4rsHnRSsvXJWsULqqKDrZ7/
kPaPdlzJ0kLZa1SiX8hGJ8Bavlt+85sQdtDu6CeL8hKHIxxJQyHMVyakju0Sm59nni3FcEAtoWvw
idiXq5GM4TNW30pVjLfS1WSUGijwGhDjg+ZuEV8KayVzmzC3aNyos/zi1gpwWb57KRsNqRqfnFn4
9qChbBeCoqTLG7mcuZeLXuzePwCNMt5jbdsHZpUzI++jpQ2hAwrqHugat9SM3X+2rtxtuoBys075
bTxwv85W3lSJ7jXUrCBXVjTBBXP0ie0lzx0tvYhktsvEjHWxeMa/of2wjqS09/qrNGDNyJKZwHOO
RxS4aoFkJhAehMUnG+4Lbl1EARmOqtu/oUZhX/RRqgNtLceu4pRblmauW0bTd4gLe5uz/lf+VUM5
Kx+s3WQo4tcFUsd6QVsDDfphSGT6lzO/DPxUdJBUKoEoKcLrNTAuIyK/Kd+uxqHqGaTl9fgmOgBg
MZgzOSa/VzqB77IfyAOfqIrl235JlOnIMFT3lWWyNkdd04KbvVcVoSJxGrQFRkTzthNBo3hCdief
O9O2EAFCRjR0dXlor2neOpEJX6TI0hZz1ybSqLcUFhnXuoVhV+XYCHsnO+sjyblJ7annYGcd0rpU
zTYfLVnC+4+PQOCCKISPVG7dl1hjq40y26tPlPWoe8vDXzy+lMRWttLCpKKGkBObFSF85E7d/UvB
dEEFjbTbh6QmyQ0ExEhrxwvN6vtXOiFo/kbqkwfkUIVv3U5gmsKHeCAyMqYe1hynmylxRGzpyQGj
tyWrw7Slf5y2YYL0+dZnwgm+i1x5l1VHmxRtccZ6VXzD9+cXAtU5cZej3fpinr0ruMmv5BzbTubM
aRCNjKXvvKqq6rBkKVbP01jgYfJCkaIkuR+fWEEJmyNbhh5Aje7CXOSpmIlz/A/qrwoF6Urh+M/7
LXyabYZji0qdaopu+dmG5xPJEqCxZR7Rtyf7OFA3u5mkiLO8Wz62/l7B5ZsGJM5d2cZA6uvIZaUj
sYZ8GDygjd7yfkWOzr8sXHWo6DWqR7uUVU3Qy2ZFaRPBGM838Zsd2r+W0DhfBBt1wFa5tKMu3SfR
cASJayeCsRTslELwjJmVHo0JhjjBccTzKlrguYZdoAgWv//K5gggDVFTGZOGUjlBb4grCVSNrIis
fT+AZ4MAI5C1KBU+aJ2MntSAdjvt3DAypBgq1+OBo0Q/9mSRFxzWW9VqcGNkvn+uLDzGVuBDM+7a
vxxcuvZ/JD75z9rpWAtMzLG78XxxNTxLJt8XJisoI3LLXwMtemUzqsE1LjSXez2540UNoF/rxoHj
fZbF0udG6Zyz0vcAGcoOJA1vD66+rPCjRh6xHCVa/zonSv+AVTj4gb/Zj38SNYbwa0E1XUj0+myz
leCbwGGPCt/Hw+fBWeDQaDW/5LWKXan7tRrHIAaQ8DGyJqKSr6vfNhDXh13nvgkl+hbXi7514jCu
BK31Of9sxeGmYEn9M+ghrSyvasZVlSh1mHcPmLI4XCrLpchC6PrkLgAp3t+GwDDPoBUsZ+c9gTXL
WpFINJSdg7OYFTRCTp4CDA/ulvK5KoLK3sgZde6Xl2lDJ/aGsxlZpuO3PpxVc0/BiRkcgegRjpKZ
5CT+jGVV/0mBhpWMjvl7+aj09nQtLW6cpQ+5vdQQ3L1uDHPcX1SxdjbCqG+kIYgGiMV/nO1bJ2WR
S18RPgTWoUnSJiR3eIDLcEmU1zhCAu06OTKVRMc1Yao5+Lm/dU2EERVlA1u8pHE5JxyEpm2LVwsI
i9ysyRXHCYAyTKvRFhXmMPtH1X7GbYeJSCLEvSCj/KzmtYwpeH6Gz53itnE6TafcZNftNeFUTU6n
xrSDLyuarGLj4Zu414mNHnjbctkxI3xb2o45Io6F9OfqkuUYGGKt/WViZdY/1F6/g93qDWsWQwt1
x6oNWvwL0HDSYk34B0kmIgEH0EY56bKTg6pAkD57ns5HfTrcO/bxmlXWV56IL3lLXKEIixgecXya
FqUwbjmve/2ep1zkSFlcuN3BCMhzvEoyuJK3AS8NddNWnSpxOFX38Qaf8SuA4GWdKEKxhjbwI5Ng
YabsFffdlPlzmpNBzqp732uG8azXWFkWKoYxxQ4MHpsfRTxnNTDjerV9KMdcdv30STJ2Kt/kEpMS
hDtnAnY8d3x8zhI9uyaTWlWlClMbob3iHJ097eoSze5Oq9eYW22ySkygjO2UJyQHRLq5Urb2jIpp
1ukgC56A7Y1khFFDIfVtbF1tofLM/xuA88CN00VC2W6nvw+cX9vZfHPEsoaao7Z3bEZz2ijpD4tE
c9o/I/CHVs1UJoEmpVNmwXv88ebbNJ/0IBNXREc5yFKYFQA6qPZamsjoD4TqVcHwpGsvr4MC2KUy
eAvhXBbvCqvDSVIYMkQtF/fDDOsRrPCVpXBMdxawAUITIY/uTG0Frk3PgqxAkxK46eFtnWjxDOTm
iIWqTLu/ygTTLl2hHJuKKfOagdAB5Sd+3WPe7McIggLILYT+bFoeyX+wyDwtOxI3P86f4iP6eTSB
KbVFc6I15nD5Hl0U3KG5OgZZ0ggIZ8EV2LsFq7c/nqtgWPBmw0KfwDcr5j54CE7yBgtinKD7oxsQ
4vMoQfLS8g2W8jSzypH8dNc431jGX9fh9gE9Ae88hY4XX/JTn6kmtcZZ034eFC64VWT/U9O85V+Y
uQpOz38DvcLVJCNEn8YJA2diBWsiRmOCj5Ce2Ce3XEK3/lCal/03HAdZLguDazv5+bKHyv5kS8qt
0teM6FVo4KNZtlnfP+WdGqHTuaTJ1YTfka7Z3X+wNcLqPt/5eE5GXAYXDSk3XzQbXN6TpoZH4uLA
YgjTOjP3bou5vU7SW1d0zDA6w9pCo31FTh8jpDhPQuRHJg0hajioNdcVLfaoXLLYzSj3FWTu4PbS
wrN/+ljD+JvVOvV8W1J8Yc8dBl9VzX5gcTPTLmOFIvLFpfEEnYs7XsAVsdlS0xX+uG7WTB1sC06h
DCfoHo+np0sUfWnbEE1klhiHlYdA5z4DPe79+SCWUWW63+6v7SgzmlhSjEMe2u3yB0YndR/osmC/
eXZacsAWC84bG/VU99o52gvMSCu4Ia9WN/XfW5jHl2C7jj8EjD/NbBSwKvREusEf55SyTwocpDrb
m5odtwjjEHHlDUOVVl8qr5NhQs0x+6Iqf5SltTSneproojzn+DTHlAnrDYplE89b8jP54MuDnUEM
/S4Ihh3S5RToUAGHyknOySIJkLvZGMPkJDGeb0u+IoeLQtYtGmTtUYw4w9+JePSxY9zi63ZcU/Kg
SZFbqKYR3evsQrOrGKd12nDq+oiwzv5BNyOC6EsBukd1C1qMSEC29b6L3INyfKeEAxG8VnG6uRed
rawWpgou+xefq/KFdzNyblxTwpvdKgMknwCrwvFwAY8fjiZGxpZqh2xMj0JOeUI58FmVPqp/oQBq
spvfAEUMP3k1/mtWquxcOndn2Cm4nLlqDhi3Zi3hTG/0j7aC/ZS/RGmrx/wBHfMAM/BGtzUci8aN
Auujl846txWSqZ7SosudzywcyQEV7tQjD2J6/1N+46/q/qMQIsRhAF3YrET0JzhEG76HqEeOLDrh
rR9Ew2je4Jo4B3cFxRi/CyLTcQjJa11ix3CnLhJC4hTi3I+30qcBv4hmzPHLXNbA7rxRaRa2IoQL
0zCiifMlbMidMabnTMAmtsWidiZAKwEc/MsdGYSUnYtRlhY8q6Xtwl4Ul0yV15qW39f3Sg1gBtgP
pZSvoi2qzA29tFGbDn9jWFX/UrITLFy2mhsMHSwxWBF5Ulfg34aI8Dfa9KpbjEVAGjWUA9E7gDSQ
gmR5GY1bGcwt4Ds8s9gCbv8q/lXB4+tUFBLIUlIRbt5DBIS1Erk+Q1OeHcgrH18FgjHmUSZAbbrS
RgDvmCrdZnoaH+OXH6afzb8EntRGx7I5UmiXpDVcV+H20Zf30FSiaVKZleoZnvwRe8mh3RU2rDmd
WU7s4HMZgahjMtwxX+RGjTuTT6Dpa7gA7gfJ5ZdHAUfzwt9TrV5W+y59OMZ+4yuWYGUsU32uhn6j
fCAxE5nWbgvyUKdko3ivFS9l8QbtQxiGMB9chso0ZGSeAGqHcriZxcKYc8Dd7OXBuOEdRKgcNq0V
ylQaPVFHQCqwu4m0NBAUerli7/FyT8jwEZs1i+TD3OiaLK1yHFyOHn2ZGB7Gr0Y6S9+4TLa0nwqy
TdPg+FIGJPXIyERciVbZ69OCh7Lp1j8yCgLtwqWBkXUxe4EHd59FIxW5d3Uwen5uW4ng5/ZhzN4g
gny1/gzGlqwBurUIv4GtwCCbp+/JjJjVB/v68iBIfNuA/+IB+Zqip/g55trgc9p4/VCb0t8GF2Px
Pi6OSRx9lGO9CGQ/QwQ/RoC7vvd4BgwbVsejGGWFH4On6TV4FbSfX9Xv9Vy7f7iORec/SM3jL2PF
+0xGn+zQYp9uhvyjYO2gqZv6HgDL325P9g5pbvmJGYMZzKM3MoI0cPw7KspzmoGNI3Woowb+5tu2
eXdKdXL3TjF38Aoti5X/jztktPoekfnzpnLL46MCN4Euub5BGIDldLPT7Yl1oN6tLBzDFcBh/2PP
SGSPyAkU4ANN9T4UtfjmkJXhMwRnv8e6u4wE849UaKw3VrQD8WTyREZNfGxhpDy4Gf/xmqd7LdMZ
wZEG4nyfsbjcE+0ZkIfekGTO6mTDcW4HO6I4lXf/73SJxgi3fLPZdiCcCcdlqq1WEAO25Jij0Htd
0naNqgKu5oyV6ILRPkOgz00T1opMavFCyy4h0ny/BgWQlahY7hAzHIIVecIzHv2SrPElQeHCaH7r
xsHYmjQRXR/xeZKQW16SmdkQOH+oRxs8EQF7AYZ8lrw/LjjB2RCFLzBU21Yga4QfyG8Rc/D7bASz
BJ0HAxAV0NvyJSeqvTDDO96Z4Ttnwia2d9jD/Qkvc3ft1nZ/PMTPGqPeYb1xHyagRZk0lKV6CLT/
ywcZ2EuIWmbU7CAP/3AYsX/Ox4MmUmbUtTYD0YkotN+LQ7j4oJtJ1kC1jJFpt6g4OLfvxlzh7kfV
6HM+BcXVdcG6JdFDAv5I/C3O78UdmM8vcg59JHtyx7kwODkbsTCI5HTMSzRASNZ9H+CmJE2UE7Ky
hZK7i60XJLrpI941LwOdfbRwf3pljh+t2jAFk9jMlhOCCOHu7vXpTB81pa9uD8w1fa7CoxZkn1Z8
54VoIVEKOxA87YHiU9wP3tWdHch9riUfrTs6/jYovVtzAxmt151vg1CNd4L/wHhuwlCpKPdORq9s
VcwJSonzZZ5rVEj+rQMKcbhqhl+Spl6ZOAlS9zDmBKpLwcAfklWyWqOv8qWLwPY4RoTCZk7L+Zmq
4aciI0hF1qBIXucrHHiwFPfHDZTt6xqo/wD9fQosxNbJhGgVvXpNgYDBho3EbZC0Cz7W8REhrpkn
c7QXjdjE/AUhAJMxowBoTJ7ePWnS2yJWONkZ6o7bxnvM0ZK8BA4TIYxNbsnX/ARtNE4oUVXD7WRb
E5QgNeLFrj/H7CuLEooIioVcUbsojOy/aVC0mt5CiryN2WK4lW+no4PHlTvdBW5gao0rqmvXl0dQ
qyPEWTGNcvD9vUo7WY2klQlxpsQp2rTEbP7HfJHljJuXsOebvlCbOLSgXGjLfvBFwZS3c0rpjWJA
RJ2vvdU/Rtz8D1T0mR0ToMS35lh0BRZJQekdBxN8MLb8y95yJQOk1nP+uEiMAzWyNCrCtyJTJmxy
1CG++pCj9lv3VBzBukIPWQ2T35KQnyEu9BZb2AXQ5XNHk6LImlY5AjQ2JuLwRMYFy+j7Fx9BElAS
4gEOI/WHnrpwg9M7UGNNIPQ14IBHCmV9OXpnXE90vBxqkEKW/cpwK/ieO5150m6tt3UwQqQgN5MC
iT5f/Nd8RUs41nhaK4tR8gTglXQPtHRWje1WnlP/DYqcsJi8AYZLMN0yf1oXnlYlwtVY+EX5XhnN
reDk/S5LkP5cnDHWBdgf3D/VrZuhKHaIKM6ZejQfCjExy1Y6LiiEvhVYKH7j05SZ9apNqvlwd21B
Rulq2a3WRpM1WZnlHQLP171HAv5HNsHEUcRYHvhmDw5fZZhkFf60WrGw0xHjpvDu3YKfWdYw5QfU
FSliaoZU5cAj7bDa7Dxw1dvN41HYi4NP1RSTJGgkTzZzAAR5jdqd6AasD5IhqnD8qWei1ndBAmpF
+VV0OCXGsMm1QAFdevCfljMDP+go9w/oyyjfu1XVGOokrBG0/FClZtnUN4oNdjKSbuyep/BtT5Nc
BPwd9zSrfhi17/roo95coXg7aFeost8Uj95FfQPD0uD4fYRVWlCs9uX1/Xh16XrpiXLF2M0mbfVC
onQh/MpmhxZI4ixwguccIYXLHndjH9yRDm5ZoZC/ucqCFyzVSaJ+wSjzMKBXQ6/9mODtZuNfRWiH
nlpeIGZaOgJlE+hz7I+zgQMvuKdLj+glsDkFQSh43cP+UBO2oQjxJMemYiXg1cj3pJsQwZG+rP+3
q+VYstdetqiTiH8QAblpB0u0RukWX8Oa2nNlRH/e3rMtxao8N4+X9DzCq71xpGdtfJegeJvcKvzG
4v0xiZQ2ZcApuC4o1mmJnbSdJG9OHrccMMyfGJrrJIWQ+lnprdHjOx7pjKnvis4w3RArHEIaS6u9
IfO5tveEA676Frr6/FJ00e8pAMChXwcC+YnT+UoUrFD0XHUeFBHoT2s9Q0jHFnAhnEo+heq2h6q8
bhVYEf+Rh19swDN56+YIUZkzYRnH7l6gUiQ4tbYTQcvpyhCXENqQnKWeTLdotrIkzOi0zMOqQqNA
S0Ckkd03vwsvlJ0prqBUttmnWpsnyxfD3gXPvwsLnk9QztBcKDS7h8k6dl5yB+lDPfUf9IGbwSAP
YWAwUzwpov3SWStQ0Df2tYaH9SV+NpszGOuTg25IynDihYoCtHIPqRrbTSGBlbwBqeE/QJP/Ambm
nbCy59oSUaVXjdV88n67iTzoRHY1qwOXJrlOw9KlZb8pdg813pTJvGgq/DIseu/Iy21Uv2gBeCbN
SEB/vOBFJzWgJamRlPzOUICErA3Ta9DZKhYPcNiss6Q9vlGxbXF1UciNdrtbBEsATnWVmAYaZJDz
cHtA5wJaAhCzJwA4tcH6L9uf80DZec9wjFLinwEjc/LDLGusY37Uadlzyw5gvlyUDp78hfOL5bLH
jMoBrdpVvOyQJR4825mns5Pc8jbRrYxfdRyVDpLlwJ8bxF7Utq6IVjBXUASMmbjFye2P9OVaGQxE
qjrjJhjsTvrMI+hYyLBy4hsz5dokrVC4wgdEI12apCz/c5QbQmYfcR5E2ar5D7drhlFIyYqTJz4t
M+yktGsoehqiDPfocKaK4lnt2tBNwuFVHMUsK1IyljWUgZfpFUWvpvdkXMN8zHPYgQrrEMwcY8Dc
xxFimBiK/ceCAIIJ0crxaRqlN0ENacLtvRrIr/aINDGva3RiZ/cR/Lo1c8BONd56PtB6EsShph1J
7TrOrb/4tii5vpxzis0c9zikDIOLlviqL7i6t7HFuQVtnjgMLJ7Gegwm6CGkNHHCePctIIPDUyjB
lxe9QWLGOSigsSEz9pqDJnxHUBNPBbnvBHx7LbkY9cP7MFs1VrRLJLjcvT5Sbwo0lv9QxXmdw2GC
FwmiuVccLvEqNusGMJ9xbatrOu32wy+tFRRQWESG0K3wuIPKU84+RBohDY0/MVdJewCN1jmhflQV
RQLPtK4zzoIppYeIEWU4kGB54umREoJtuqF/3MfwEu97gfIqfM2+3eb77gcWa/ggCK0O/5G4CszU
N6owRlYusZQO0RNht/ysBUF4t+iIv16NtoFQGKfyBq3AqOSpRJz60RJbQdKtMDWoSqA3loYYzPmr
IvnY0xCrxqp1DpwF12uxM9caLzD/eufnrRmDrT4FEoUrvzFMJ5kuXBCWJwdDFfkt7fEmpNyZCdK0
x1EQrbyYXDCxZvBraxcvmwoK4gNSGWLNjKNoyDGt2VckpI49WD+tzbIcb1e/hZavZLYzeQ/rcBEw
iMAv1NLYOJ1O63QUV4rjqA7LhxrdztZArJZHW4+3pCkE9OaCDSSYsNXjDJU7ur0E8MeCicAbL6T2
ZrXXFoIa3Y8lx5A0uibqu2ZPOeaQjiVchdDvtV07XAOtmrFIjgmezjOFN0I1bCMbx3bJpz0JGjcr
8NW63jBHOqjNzG2IGQ0lARnOlnABUrMDJpZtRpevaLY5wjAUmKVyxf0MPRArXf+b7bW77X9nGG7y
Q+pEOmUws9QaHK87hslxJwIcnIcF1qHnQqCNmKX7shb1QwDIuaxSSf1b5u3DrE5YTgWImHxIv5ut
BjVioQlR6rMYUZmAdkRd4lQE3HqI8EmQXF1aFXAftkKe1S3was/bmswjBgGJVpcNN82O0QI3TQQT
/0RoMHYNE0TMV9Or0dvKGMgQsps4F8pDF/Zu/EjHrDkqnWFqy9sVLG8Y47dHMmMjc9r4yLEPtcE3
/p7dSIrP/K/rX/TQy65kgpUND2DHF6YbyugJI94KtJYImFN/6SIObzCScyd5fkmr/SuBb0qcLTJM
7yO/IwkhI5Cssj3Bm6SA9Rn5l8QyuzEnOgj0Gh0sb4rc+LUNxpguoyx+Rdbe44E5j9Lm55UTOkhm
HQBf7gxrr0NuszlAfIBibo32Hkqebvye8imBIE9grNqbWO2qq1hbx/FMj18PGTN5KYOeMPKQ3yvk
HnXbjmvw7hu4anYvhfQ1BrYMMT7LyfLm4IKBHT770WlOLz+G1/Idm9GNWr9RO4Jx1NnKbr2irIFd
/j8ILHbHeNAKMMTY9VFCOPNLy8MrY/S5VMn8AYtEjk+jdqUBh6TLhRC6eAAKbgw/bMagiw9LO88S
4T+CJoCaH7bI0qkL4XD8nqPC9lUWCjZGTxIIEXAvVzI1eKwU96UV0vITOx5uny+QZ5ASV4p/dhPr
qGcwsNsClsDjKB7y7XuVW5Q/nylzfp7SsQLqbAS8nw2r3YWAo4e8vwE/5XJer1SmWn5DP5gxvLib
bpvrkioU25lmOJ6y4ZJy6jVNND+Zpq5hy3f+S6WQ8LWpZn6Gkau+fzfpsKXDup+t/dWEGJOsOhKv
g1DCr8WhwM98Sti4CJr30+wIOApWv/JaOFidJ4ZyKx27RTyl9fOOQyC6g6rWO/iJguESFLBIjKFY
XgQ3dTpxtoqQVzVPjsc60dgMpCrUK4Hbrru+wlDvLzWOQ0HB39l+Ox4N6QV6HyQdqu/VbcPpp4bu
Kaj0AZ9HZRsi5zWeIIl52ICnLaGmchp0GH2YoFelFjgAllhZVEzJ48IrxlolEdFPcCGgWyjOT4tD
hJ+5WSF7GfMJaNRrNKicOUraBQS8c9SHMGjxWU8jO+nkH71fjraexIo9vwgo1kBwP3/pxFxdYhdI
Rs1SgKbNuX+izhIvYrTOnFvndObGIKFVv9uw/JUiP27Kv9Tti+HDcO6EP6Br1X2c3jPoqsoOBdE2
KeIZWgdpYbEtGaGKVWqOIx+OscDIpuK52UdfPqJpNspXUWgPOPJb3sFRtdAAEXO0ef2flU47qJbm
sNZRLi1q7T1cIo57CpM+KTDAeN82HI9zsT/dlWPHlmn3D1wjmzc1qIISC3b60g/XLFBPblIwTiy7
XtX2YQDtNB2s37JSJ8hN8HlFBRTcHno8z5nL5L7OF6/dWC9D4JASPofCZxbu756O5xWB1n7lMH7Q
ck4enTEFjTmyufb4sIr8/UMtN/0eO9Q/cEqqkVCaG6rwNqZY0RuOf61ABxBEf5JcgDRzfmQFhIyP
poU0jO/Tzz7PX1aAdcTNBiCWCCIxpDN45LdKdFHvW0saj3Q+3xiNJNri9aAiUHu5iZX6A7hcU7L0
KPrjInHpXZU2rgCrFtD9UpiJybFCpLWHWAfm+HnbSSuqttFMKGmjWN/c1KK8H5Yqvr2DhLa+9s9c
719bLsRPc3QbmSSCgFzU8dqM0WT8vshzd4pgl/vWomGDF5eV6scjl5sHID2KyMsJJV7znZorbEkG
gc30AZuO/WN5h9YvZPrnp1aC0HNAZjYu6keM34aHyzcC2z7frSKUIpZS83jHCOR6lgqqQMkCTZMp
1qA4B1G9NTtnjmnlJ6RXCUDx56NB0pZLiGzuOlAorHNlX5VfaWOfqWG7s2aQcmuqWrYyweSKyY1k
21XTP26Yk26GxpfdHYd/4+mNEtyUzcIWa/jDrabNkLQZ8QjLHXJ3f9RTLzthSLGOHiTQnvEivUPi
AHB2XOSkdxQKlly4L2eOsWVZljkjxb0jpRVBHG3eCVdklG7n9N/tNEr+QCEuLisHVqW0Bd6vVP3H
M0lALI5LTAG3om1td8zhYu30TPfTLqNRAV5nr6yizqoWlYmwdwG6kudGxumQH01sTvVPY9mzZwID
c9nt/1MePhgvc6hMoVA0AHxa5Y1muHr5M7hF0hpg7AiWrI6tHJnK1/lpgkeolTapvh1WoxOAou+Y
GmTCV9ojbDKREQbNXAIcZjn1sz+O6YSsAEXB95pDtPe+SXAFNM54bRbwfDIm+3c4THoTSTVc7Gmo
uv8Z3bk4vIRPZFpMTRzxSrUmPmZmmyJ/55Sz+QdYKMA60bjqppcgrZ41jnivontNxq3k/XWHSNRF
0/sltANr269J5gOO15R4XjIlP3u4CTeegjz+Eo1x/WA+JsM9G45FAoHXXqVv6Rkygb8ATBpqs3Vh
uTTaQ5cGOg/uWU5FrZi5ARKqc+icesRaa9t7l1gTHzu3k1tCvyhGaL9I6d1lwfOQO9OhvuxqniD1
bVG3M8VJbSgLiTkDM8NFUsA3vHjwMgliFCPR4uYSGXjv1VV5jNWWNCPCRXIqQcoykcsj25ZBMiOp
0342haTf8amX5xuzvStB05QvVeMe6KqdMOm3nnSPrOlErlbP+AZR0qgim7FTXKutw3lh3YcfQBOV
3np6FwPmuuJ8OwdkRxR8iDNMK1/a4JploeROe/Hw34hcgf8/cFAmF3q06A5Ex+gn2n/YOD7zk3ul
DyAfz1OSlFMKqtg8/OtX1WqvXiRwAc/pEzIvAgtHXw+utXY1ZHuYN60Z7pVbauqBFStE6nUTee0B
FN/MsbYZ/VPktGje3g2x/qRnVIIuLdZzPn5uj4+w1PpSUD5//jkX5oDY5d4Ki9YylwDwnB1QR81n
EcxvNaRGASOv9x9WuZ3o8fg9TLJyYZpDx3ubqTVA+7ZrSXIjdPhHZSTxrrYgar1m5uel0LZtCSzl
NOJfbvhiq7PWQJ3VJxM0QgZWLdezRBGT1wA7+kVLtf/fH2Zpy/QR4zpmE2h0QiRMNwu7SMhyMXSy
pPfxNAP3R78nWJEy5jDwcvBFN725RT9tsUzXDPpiVtk2pEie9J5Uq5FicHxp2tRz7qHLSZlEgS6E
YLOQvG143JhGqV64IY55QOJIE6I4Ucw+b/pF+EmJyBIRstut1IG5pF8tDem39/TcwNiPcQoc6Nfq
g/btDPjlFdkvxlqiUX3bT6dwMhJ3Naolu68SRzB1+eMxEhWvGX10s4AuM76bK2QsarWFvB8mePF0
7mZnh4YXT2XV5lrLNdx1HwacwoeAEvxlC8f+tWsHxE4r7jUJxEZU313vmiQD02+JH2jxIpTyr9HL
hgEHzuA06oISRSe0KYmVYYPMIW/+kRoV2kt9rdU/LNW+gHj7Q4aB21I5LGWLwOpML9kzlVFMVWJf
4lqlOIY+r872VtYRKuf2sbk74FKXpKL8soc4m7L0yw9nEMyxu5lt/NpP3CTrEP+EHljNfcAD+lPv
qIpmyx3DPZsAI7nEqaQGyCdDUG/5UAHO2HLAt9mV3O3w463Dcn5fw12ijmjyEL12fD/4I17QI+Jc
EaqaDrdAm61FYudt1VAgnuBdd8cF5134lWqjM6hLtsJRWRJAr8KMfD/bWIF6pvSwiHLBsYfybbmH
WKqbx1F3elxfmEfqA23clTmehvEcs16MYvNoi3BoRyo+fXa/mZ7nZeLx0k8h5B/ANswaWfF5Kydw
TSL6OQpQBaoJcnOZNq58dxgTEHiWa77JhyF/Sl5hT3a4QNmscMctGFRk8n4z3VeYv7WzVkh9tSJi
L1FPxYovh16uwHOYzhnOPmqYmXvr/r6T1gPBCnBuRExGC6MXKQMQfnoN+34T6HQGNGgcROWKmZWv
iEF+cjDygzZ0H+QS2Yt0LFt1qz6yoiXWuxVIOSSCiqxK5JhtPbZPMp4kP0a7/55JsARWPW3fxhQU
cFyr+3RANIMC+Esb9vq37kbE2fclTrZJpbo1EmqB60Brs8dWjBZTCypZfAuPKc9g+Qk0nZhCrah+
E38PUf/PPQTVZEQcYjRxV6LBkwjdro7705etPOZj1250SEi8BtrHKBW+ymeLm/H0UFZIfWjrNgQi
y4ZajXqna/N0EYKFzlkiiP+IWCZK5RWezSvEBQZx4PXhA/afxsP2CqYa8yA5JdcVGMvs7IKuH93a
MFvCsfy3boDIDkkT9q2dAG3CuKVWzKp9TiVesfNm5bxIUNYAJRlvIGUVJwuPTVCbDo9UqOSUJZuI
mZ3P/AUfT2tsxh4mKk0OG58Pu/1LPYpPLVkS2LzITrNT4zvH/bTDkOkmaoAFAwlVhAJxLGjrWFA3
0JuCaP8ixrP4UKUHmpPAQO341ugRfyMJf3yt3E4uItX7uEAYvk6vpQp3Bz54eBJi8R4oy9pXtdqf
gxf7pS0KjKizFrR6Xw4HxZ4Vk3uk9p5NXqbFLEjhfnX0VlQcJALItYo4yy9NW+X+KxHdQ1yKPaSi
BJmkwZB+gRA7vdEn1JmygE/aCJHlNZB500BqJe27uk+BeZka6cQ9bisV9ft2qY6TGBSKu0/3B5R/
pEfHGPMTy/joPxfK+3Aa4jpYSllHoe4SySjwoV32KX3YYJo8g/CI4uKHj9RGCGXnrOND2b2E6o9/
IW/fj2qJQJyctHjSdheHvJuqHLvkkfDV5ky/IR6PSIqNbxGk5jvLmlhCcwDu0AZxjKtDlst+qxsI
4nwmmpU9XqVQIRV99pLnYDC0k+OGL2nyYozr5m77CPN8hfGEdMUzzTkqHMu1b61M7BotCuPf/YCi
1kg2FDGwAroluxKjU4d8UNFJ/DSxPtlllat474/ubfJIdpju4Ij7Ar1cka7AfyKfABLBGwrsvWp0
8jqAMn+ZM1Hbys1BpbUv9ciKKYrOVhlVbBSchXOru4K9ojFwwcZjn6A+6+uj4OkrNgoJwEu1b6kD
kYGZxLv7cVZ77zrq0CIg436kFXj/6Q4MIss3IDZ8BGA6OpOIBqDpI4GP2Dcdj6Kf4ayLuaHpcqnO
KTgFkpolPFVFaIOSYc4viHqz9rtznAaIk/Q+NZx4iHageWJFpqDnXW5tpuzh41ggsVDnLQg0Vs60
PytM+CubK4/1HG953Xh5FQ/wOh5y53NHXko+M/ilfl2qeXENtnLCO5d1EiURjymgGXDCCUS91YIm
sx5rURxlei7MAqsw2XiQ/4fukzdJESbI6J7yrBClevDWG1x+d9NEFzMRKnS7JKEW1/Drun0G7q30
fbZiUeq47u6XGmLjsvk97m0GGUWtHeXGx87BcS37vC3aMn8XWTM8Q89VAw5Qk8jbFbuV5Ttlzr8u
smZgwHuB+pF8HzHBRAuYBCzWnuOUGVMgdes65h0G0LCEnEmyayYwd5/ol0UTBsrljNFclHFXahcR
IB8J794qePde6HcQ6Or8AicsWfxybfENRamlta08htoliFTf5Ccwv6iY3uzTzm8RmnYlMdsrJ+Ql
sH82K2FkdikOTRhihsnKmOG5viFqLWB85gJ75LX9+sRs4i9bW+TGaOeqUoN0TRH+nZY5UHI7kv46
nh8gdPiU3vtSkX9eHCiIaurqlWmvToGLp+g3pKtWwjZJa37mJ3Ge0aGRVc7d2A6VNMCB0abSjapC
wQ0Vf2paV9gbCn2lyXebtAHLb28kZwVpG7WsBL6tKJvKmLtap8zmK/sF60wTX+SfLXhO2tdstjj0
i5fUQ7vdcrfSFG+pSV6nWCxAZVbvMPizQVMrLwxhgR5xJWzZ2easuoAk+UH1KlcGX0Ua/YNB6r2W
f+UullvBwQ5lHVv27R26dQEOQGdK3oRf/reuc5nrHdAVlqF2WWoakz7iYQCyvE9OHGNR5BZJVeqA
oOJyEvNAkBqZqCjADs9nUnLMAzYBNRiz7wimMFyVE7Btj2EUMfrko6A10EQ1AquKG2lS7KN3dNYK
gAgL+JXTg/jZYPoPpviRCkRuhUf/Ulq/Qo2mdSgTH+W51/w3Ux4ON8pHnwPZ7nCcgoyZpg+HkJl5
bzMg9Ieo0P2JsMrRjDZsb4N4ZisnLc3XcmuMNa3kVzkdaaJNqc8vbz/qbjXiP+8muzMliaT7WYij
o/9ofRFDHozBwVHm1zLjEg/xwpJommh0sbWVu9fZivtV2q86Juw1fMP7G3zRoFXHfTYKKydQtZX1
Q48RXhLj/tu+FQ7gejmYSnY8hfA+1x4WmS0YiIS0FW3Xy/D5n0y6YrJ/T/ISka4B0xn7vDra+3eH
SrGQm6IlW1z/6khqqvU69/ee5XH3rxkKoleeEC7Lhl8eM/5F3ft8oPv53RFh0Q1Ei7Tw5k5ubATP
nIBDE8irmjqTjN7yfP4sfNFEcEvS/8d82W+slrYKA+C03Lg9hAOnCRc/1i778XVk9Eu6coqRK9cM
DK2Ck1/9qsJaozJS2VJIz9phcKXyAIw5IRHFIWePe84X4b4219niOFqskA6GjRU0mFGgWjhDIAol
P9eGvi7fWOpRcNDpqZGtyKYJtN5SRCQzF4woufMBkR5lzRSdk1d3CbsH90moJVHvu1NWwtQcrdIX
OnpJ38yt7YN99e5L0X2ViaWVYaYv1jU2SNZPb2zF1Ta4dTpT+9tYAi3Z7ATPAr6HZMOIf4rKteIr
I4YXbdXLZ8wS8MqWUvrp+N3q4L7gwPhwO4KbivCqxSccGJg/Cgl5Sag4yGHKyrr0O8RN13dCpoJv
Se8C4Zbp4SxmdiwiN+MP0EZfH9nUkhA6yQIz3wvNg+Y67MiCUGqbOcCj4wsDLubCmTvglQRCISGL
xe84TRMpwGgppDqtDWP1tc8dX9aiUEP4uw+jwRhud2DyJPfCqWGTjRupgOX9Bz/bAnr0ViSqEdxL
WmLH3auO0HbhR7CSr4zQLHntZdSPnty4DAeGKUu4ieIdOjilrnRNmaQwnqJDnqqg0fJK+KZCF4YA
MLKCQmwBwQ2yi/cnbGkqjr0O/82Qzsgb7weJmwKbQLCtjIdUVnNTklaG8qVgThbsxenp2ddpXNRL
hKVJBfv+VGBRVqfE7GgIwgHLshtM5xJ4u4mfvFkrrPuxHuibNxAWTMF4j9HxgmRbWHw5pFzs6FDf
PbaE9Dmz1rYmCfk+FUp8DivzfKQD99OMQe6S1HzHiPZyVkdX4+NczrvlM9I4w5CF0okqVgG9LpYU
JYCIwbRXbnErRoe3IQn8wqcVolLvsiOTk3yCp6RdBvs9RdyntenrrXZidmO/TaS7kqCn2D54EZ1x
LhaIemcKdhcnA1BRe0gFeLy491LsT3DT9c9KGxUo3pGITr/y9crYTWocDvWJfoIg5FZkV2HlPTox
SkXnafYgIPWIXd20M5Zqmr57lgg6+9TRQY67+qmN83n9Q/ilBUMmbQcGu8+7wfIkoLGvyYutMWoA
Jv7023DGTJZtRQ1be3GIHYbhmbqpajYLXm+GUtaafyQGKmpzoWB6MXqhUebjj0IU0+/5BGENyaPb
h/vhiNXCXFLQ5LxulMMVAjVm8GE+/w6Vuf7nHwKFIF8a4sCqprwg64nAl0q6pk+JvydHpy7TY1Bi
QOGXKeo9LGJGMpvKNneDd0dHgQjiXgxAptoLcF9MrhRnbh7KXiM4KtUShAqIJ7XTj64pRU4rDFqL
zLI0BhGWu4FWhxRGeJ3rsebaXtLvq4BWGlj4zo7GCgZ02YLowbiYlhZeIlwe2muwVhHfyrkVBI1o
gdNm6pR3sgkuCHawt6705j/dwoEjq8TAcB/e7pmdkzMOOuwstjwOZCTVtPfjsXLdNFtjILR9ryDp
40CyL/rwy/Fyz/HEz59xatWPliTlenNVKPfmNUg0rtXXof6+fgBY0qFteBZ09cwoN2BKrmoC4yuW
LEaJSjnl0ySn7rtAhJxjlKdjx9ElYtqqyIhyPaAnzFUq6q+Atpuus8Z8444mWi4lEBnC37awjxUA
D8eo+R8vUrgEUdKvpP4mUYzl8LexWKsHwJ27QtNZ/NplnhNwd1YgIbxfZl2Xhz8PFZIiXHc+hQwS
t68kpMvrzV2anGn6eI3dkEOgiY2zcn6YNJngHapCIyewHE6bkZRviQh/gB0vW71BOLJjbQ2ANqFS
r9Dh2BUO9SmrwYlifDFzS4kkw0D6vORd/j8l4KekDZYwIb/kvVyzlH8zy9JQCYFGXhxsnWnd/Veo
vgnS+ETxSUysYArgl1xkIOY6qlvkWU2L5lD7JxrV9zXnnjHjqU2AW1MeCkH3sz++N+wO5Rlq8ayw
t+pAuxgsqkMopcY7Czxhs/XnEMgxjjY11w7MeEn/n1rdcl43WT0uzTeQCrEP97Cs0oS+rx6tqF8W
eCKNQwJnQkMT1hMbxnCHiWH3967Y4lO4QSQ6yAhdXXOliljlnqR8S05ln3Y/8bVfA8sahWljjBSx
0O4DRF6Xwu9YC4JwJJCenwBKmiym4BcbHNP+1T/FF19jENsXLMZYgiurVUQlRJuAKTTLFdmevG6t
/6mJ4b5pol0qoF2D1cumo8VUNEq3hbr4SspQ/Y0vkYQAeGmD8USkE9HX6v3VRRit7yMD4NrhFiZB
yycyzvvfysKDF3bhYn2/OIyRl0qL47EYxB6gToEbRorkwijgatTLb6GuiivedUtp7jYBtjUJTWEw
Lx2VTW1Ak9lGo2sq+W4wSFixkp5pMHvPUOZLhnqi8BfpuUQeNEs8L0ggJ+zJk9yTJDqqPbpXSZnp
tTSNz1jTG8/RiG1QWz+ykAxPgZCxZde+L4i7LNjy7UW2IN7mJzrrP/oiLJOo1dwDfwHiAcpCTjHD
tc9TyR3209w3wI5ZpsEvs8LKTZmDQUuWyK5WfNicZ++m7Yp72yRvCaYDg403djc/vC/mOgxDnXfE
mLPb4eUtGUU7P98ykGUytv0C7movMC3q5RU8I6DGYlNe0K/FANdh0d31nrn/CkzoYNoYfBmP1ygb
zgZXYUsK0oHmNISm1bD7Snn0qgi17p++hhScZZfn+z4QUacdl54MF/nONcA9I0Tp9mC19JXBB9fz
o21DxrEMj512zjQGaGqNFDidswJccdOYaLa7yy6fdJpF8JAxTbd4M5C9vSwaFZgPKJlMoAuVsV3s
R89ZZqXDoNTrv9ZoIJANVnfTJwjuSFFVmbHPMGTSl8A5wXtmS/v8PUirFu0KFe5T7S6YOezUWClW
eZ32xSeMjhwe3a/pj/IKTD+Z2MNe2iW6//WZ6XgUEbcwgXyJzA6kpXvR9zP+RmoGf3M1KfEKgtae
WzJkT8cuA070rjPlJoLGgxPJFKUfaiJfvHG5F4dMAuHI/iHvCrGgZF993v1UE5SCtTU7/VEHvInB
tfgkGvkhaWfgLav8tOWpEFWUQEv70YOsdtUuduOCAyacvVzKdKbfVm7fkB27Qrnb1p3rlCEpSMhZ
dvJlYlOCEqSVlQeNJovaXIDanJ/yacVFSUqrL8gjnEXKDooJ0stwHE61mg6xe8T7/XmAOoLoOZSE
QS4w2Z+4Y2U/V8OietdOi7HZKKDxJLV/eCp4DeyQVuCAyZBsmtLuwNRhXsEowbPWxZB8dKY6UAa/
hU3EiOOb9O/6mhEhtfEL19hpUzL1cyDqRr/EtDjFeyJJYuaqhSU0BC6p45JbA/GSV5Mqxmd2/n4v
dtw7LFdxW6wycrhJvvWuKmHtSIIbI6voMuhI2AbRNUJ263t0xaXEcHl0M6nNuSln9Ebs65NgspNQ
ra6yp/m3RgejJiZ7185jaosK77oaAGg63YL8LTP8k86KqqBFgt5GxmbbyFTskOKM0PU+zPNN/JUU
Ah8CfR8GSIk4ND1H6BFnh3ulXrWfs7+0Hoo7aWGyYln+4S2DxKyp9sJmvuRXARDkHIQvlK/kQKh+
udEyz2PhQkznTzYaXF20VuloRrazpSb+f7hilH8TB4YiBHttPQ7CBxIUAO+epGjENffn1Z1XJ6iU
BHBWrroM1g8P3mKjKkTAh4Dd8MmsA0fgmKw4s0l8KQC9a19fN1zH0eIVVyh4B63RJxd4v+LnA6Lh
y7+mBv4vQn5ZCOkzeQQNudvmMNVBWBXjNWYmRkaq0ThXULAocAK/ZlldXkEEhtgL+qnyeMw0paaj
EyNaA2JvVbm5K/GwCLg8d8G5cvzQQRjAkQP7oEgHfspQUAk1Zx5J4D5TQMnYmgKzgPEDsgbZZMri
UxsIldkjDCVaC3aDlGgPQx3gF4GxOA++94SM/LEXukzQ3xOdLkdsJWwQvwqnGSEvhTfUwQIadmuO
Ih5+dgkA/bieXQRRiZ5jjqc7kwIMpncaYLkiHDinNa7Iw5QHvtv6do4sslzz8P8e98iRIDYRrPkI
swJN8+r3Q0FrmLFq7jEgnQSigm5vFiYN3+04OMvr0cmIO+2wduhCLVqm+tLYzHpQgtH6buLA+HiH
eO6Wa36zMrC68xQgV1vydgIvGEpQ5MGBtPaH0e7QTs2o+79oqQ3EhjxwuD7RLIoVKWenmKF6PUYP
FtXq7Pae/U2N85vYEBAWUV08fQjCK6LUjDeS0tuGVJrTCEomBE/GGEsZ+lQaIgU7NMMwSSIJOq+k
8GQmLEGQpP0CCejrJ12QBdCBG9YWfWhZC+d93xeMS5loX9queysLPq1aoJhGsXfoda1axea4S9KI
12BbxmXoxuXOwT1iB5BfOr1o2cjkgPIEqPf9VbxGM31kJAGWo571J4XovJ4BSiIe89bfpk3c+FJJ
e27+fvqnHDsBFJ2YkDifLLn4C78ZCNGcY9CAdWAgh2R4Kl/cHEkj8+M868ut6YucnpS4msyIhg9C
sVCOkiJx9USNtcCDPS3PqRji7piSLuESN3FEtRi/nkh5XRYr2EnnKQcMg08dFhurwa6/+DffwmNo
y1pnpumKTnjN/WoKwqHnwRseJ/8FsTr3dRca5JVhQsOQsobz7cwo6kZROUWJgmgIObfmPIWhIFwG
GUSvpm4m7rC7ORRTIVD5sFUVlVCpPBc8FG02CZxrSkdOB04aN4PjCLSdh6cHSOWAJbisX52DEt/W
cys0jxLmbAK6ZIFRr/RmGf+Iw0Selq4MjAghv18lJF7Xr2rxrLQs0pUmiZZp2xhAQFk90YPb8Mzn
CFhPVRT2vIYAHUx+uJKflXi3120RACXxwYmV/yC1W5nnYsXIe6O5lcxU5JiJIwHYkRi5eAxQycgc
xgUgkcvTB31vvLj0yo3rx3s5+ukSBGPRQ+0QOx8fIb0/ypGI+PND+tIRS05vgiFbG2CdSN0GdFG4
w/nHvWYxtqDzxrnmmzuruN6sZGyV0kHQqQg8/pI2ElOw9VOBMfZZzxul59d5cClulYfBgv9g/z41
m3waoPvAF7A5fyiuBnJp9Xc8WQNMGWWlfy8/EsILDax4OVsb0vcW3f/N4ubmCEnLcnQZlB1EXbyO
q+Vz7eG7U4AyNZmrfden+/dQF1Oj4AxOkZxavFWbFiljjW8kDDaQu+nknlg4qS93hhiRMHCDRD5+
exvbSSQqMCUOeqWAP1nMDT9ErItYLkclKlwQNRwCWdBC4PHXicJT9BYsGqDNE9alnLo4PtUF0xYo
VS86HHKIVhDw+MNX0GcPSsmJMCxRTtRp2iMnmTrJnPNmCXZ0BpPRusxpu3qsQ47TmuDu/5qZ7hwW
XwcCjNii5vWK440AegsKhHeG1RHmTwopbs2qFObmjpUAChd3qqWcFkfqaLIrKcLkdVmehVeWv14f
J7S38HiCP7yuZ3Uo7LrvUc5pVyfnzsxJB9IV47WOgyrhTgXSLszs6U6Fpi6t/WQj4cmgE3ZWTHEN
H7lC2is5GugdkA1NFhRkZL1BUMhyoLVLUviHRceCYHlzBjXdRIBGC/KIytQSk2qEtgtPDdK5ppXe
MsPMzVm5nAXsTi8gyEOLEcJ5nCsp0jM+ytLDOkV2yXro2mRN99nIKpgfmlJtsg3KxQTffV/r1Elj
IxMie0EOiGgEb5X8gOh+wppswKTVd4XofNdOAx2Jsyfaph3GiT4eY1swWCTThjvWL4/MZ5s4m44A
heW/8cEiOLeYIq1cOh11PI8gqr3cyzZD6wratDK43VbqBuls8EEr7LqW8f3deZe6f2NGp1R0yDgr
MGLb1BiSeoEXk7oTdijjEgbUZfWMb1jjnY1HVk1ZDTgF+nYkqB6KR20opzeSxWeHDtQ4W+PMcmvY
S4x6MeQ9S82mSRQskDXelxaJJ8f6vdyg90l/sFETEHmfPR8AqSBXmLGKCjEdbG8B/yCmmAqBGDNi
OqtsWHdxp007HxpH7zJxyznPWafGZj0sHreo1c/IUMoP4WkYn3H7YvNLw1cv9DoIgfhJxqpwUmHp
ihngOKFfEMXy1HQ9zPD42knb28as2XFNqvWTovd2/c4aQJcZ2vdEhttJti4xFB7GiwSsOzaqnnpz
UB6Kx9flB13UXnoSqbSbpyYZ67DCRZnSdMIp4lE4tAYYnG1LBHN7wO5JiGg9phSmvggEUH7Wgj7Y
Mu+n8Kxh9PkgSfIr7Wa+KYScZQENl9CDE0Shsi1w5og6cxK99DSvTizQrwe+IgMA3Hft03WS+mpV
btsO7ffA81LE34KSfxgc4tMZLKaWWQO4FhcQve4sTPEmqfz0R5zcPLToNiC+86NgWKi1DWkJ94Dz
XjzaFBuwYrORUan37jdLgJ48/r0SzN5KBlwLHXZ9MN7Pv/ohUxRW2Jh7R9YlhY7CH9EqpynJuFJ6
/ohngoW7yhf+qDPevVrrWJ7e7j3EIgFeGKJJlGH3oVxgP0y5J8P+vmvLeD75FWXPC2/yy7rBbyWg
969/GUQd0XMXm37MM4xyqbsi+TKWCasXBD/QNihgOuP86suPwtxX6WnRd4hZmlkzXPMDqW5TjpcS
KQI1MGH8Pf5jcnChaj3ifdl1yzF3zetupIYRG4fkrcQBAoy0jqE8JP3X1C3j8/zq0pExhQwJ3N7s
HhU3+/uHEWrN0gpBuVyEYas8nZLgOL32lfuB/bLP2LeFwdRMWqMHxwnCj36W0r7Oz8MrsYZhi8LJ
enCk9Z9Eej650nU2zDt/2Hv2D9+8BFqRKFoeYv2uHxcIm1gpM8k2/emgXcTu96HeblnhpSX0tAHN
PYisN8QoCgr2Mwhvkney+R9Tw9x6CckuHD5sY/3ZH6yaMzF1EVDKyv0YbdPpuKaHIm9HG+sidlkt
b8ukRfzqPGPQYu6pSj4Tq5QfhHGNn3xbjQ9zV9KxjKuazkmcW9jlvs527fyJSpCaw4BiPIEJI8bx
EN62FlUd01j2g5q0NhARjHVz70zouPG51Cuknvfa6X5KaLxpJJ7+VM04tObKL2uEvQRXPh/bXxT7
fWY9BLdGhTcfVJkHWAbMVN4P0OrbBrqtbsVdNX88Dom1PgNKxCwYU/8lEeyBcYuTOQckOphJiyBS
LE5Gs493Ta6xeFzPi2nzXrkqL3s30C1SxLGcPiBWfbqqUc1GayFl5ddo8p+Ib0vT1OuSfzKcQiqa
RfRsMnie2o2xZAMCFQjCZFBsiIT4oHbVQiXAILWcas6gxEe4ettTDDTPTHJL6hpfdT1z5wBk3upj
yOyaUmUqgHFqBPrxlRZLkm7oL0yELyOq3ih86Bgi9DmucftgbTzwKRY0ldWiJNWsgDfJL5znWRMa
Mx5EibEtgbch5LaE3+2zCfryxTjuMUyZMWPMoRCXbq7+Ux5xAP1mKJySqVAS0Xef4njc1NfwrJXc
SEN9jD6Cka+PZ0tq7pygflQZtn5dl81+JhaK+DZeSG/s5PUKt13sCjmq5jR65Uf1pq35hUbsxUsg
u0pyOSoBV+R8OTq4O6iWlosnHeJ/m1RJKxYsNLRKZ3Z4h4CFhKZLT8XPkcanJd23L+lwgHYh7Gef
wrHjKD6oSXmOdgJbuxQzK1rE+64ZHlBnhhf+AjUcUuHuevy+k+ULpCkfPmBOUJANeL0snuES5Sk4
mZzQWw4Tn5zLNZzVKO6agm+TPz1gnWIbzgQ3CBwhsSYbJJysmCZykCYPTWHBfjmeta4voFFISJ5T
trchpt3EIcOpVNptvhek1rGpUj6tfRyG6MrRxYhW8XI6Sem5375E2PzvoTaZYb1zwqYESsXex20J
Yaynpv093ymglNX3pOuNwj3EKA9tZpKmwDdgDfvbPE4zKXEuZ3x3wjGpVRvlS+/1GtOtG41PKQPE
vHf58YhuHpG5MS0f/QMjh6MneTKLRd7jevamBHx/fWF1L/sXo77aEVw/4gysGKefsiTOt0XQzPFw
VXdGynEkfs2gCXx/aIFLSvAlJnvjjGEHspkBC/0fHQ7nyeDYccU5WDYSP/3/9ffheF/H/JSP1TUu
zq6ObraJBh3kwptepkwI4hDyraltz3nLd2Xez6bJ+CI0OF7c74Lc9e8imA1/DTzO/HjeQ57+v4dy
xwdq9iWz2udK3iWcclhmRMykyy5anCOQn6QhBiLwoAgoCK2AUtTmDSnRByoW0yHu4E7Gq+duVXCI
S+C1oTpauHA/bKJjXmdQdFVnSdtwVqvRiq0/A1Xxi5dr3eZNDEtN0oVQ/lceWPQT5fPP89T0zvrl
fHQMyHtx+jzOp5tClY9Xgx7U9pOUuU+zoNPYFBmmjZdR54I9n5TUVcuEBbfAXYhcbnMektQtPlR/
Jrb5cNCzMosaof0u09BM78lng1+lf4LQLYe7JJKrbFbD9h4lzdDCJfxzuK0Z4gU56Txwwaa1/heZ
1AhL3/+ZJKDoy99M0vdNw4EqAlXPHh6iB0FCwGJCmBN8CT3VVi8/+DDuy/4xtw5ucBAF34nWgQ+X
WdMbTgEXUh044kktzTQUJwbByV5jkqm8LjiM+6S0BbmuVWZqs3EkJX04koboGjR1LJJAvmT5TsjG
33nwYytwBx8D4YxXPlt3zdyV9WX7+713t/vXkRaU0AjISe73b5xf1woIe4VuzRKmc7rh16YviXFX
tX1pdQg70QFEQcZ1YD4Hd4uFYougcSzn4+LqF7XGac2SaZzEcdW/Bpwnneu2x8L6KqYoW6soJjwD
807QySwkf5ew+6eV+uV9Nh08IJF9xuyfAyGlpKiq3LqmaCoKixvciz+9ahzKyglnCHKn25go0eXV
Idv1BwkQTvZovdpylbXY6FXvXdxBDp+QK+w/iG/8GsY1zG/b7Z6YOXW+wED8sO1gpvAw+C3y+/Hb
l52U8EmcBwSQasSVtJ96hOMjSz29rIcWYBHkerpYPeYbkkqayAM5lzyZivCHcgMgLC9nSEUQX4QJ
P8fVgKve6OOqcusDJkOw64/54wPAxnUWo/jmesq0pEj5D91IEDaUlKoXshEgS8o7EjeYbUoVfd7C
8AmfeX5ToJA6uDrjq7sxu94STL36DL1GY3VpF7KwUTRQYZtXANlhKjyW1y6Qvj9+dS2kfVTUrRiX
r9ywh8N84W/+UFht79unzDAwEMHCU4pspvmt9dPFiSic/2NQw1IugvvwnINUmOxADtLou4XcQ8KE
t6pzE0lOGeViDOrIxfd491oSO0bsxvpTfBuFvNrovgXZeixj44fHcSGG+/gBlvILT0jRjDOVgVSt
VAXqbVWxOFVFIsmLPlFGLiKSlVTGQxShZJyDvsb+h+6AXfI4hU1cMZh520j284n03gXnlvSl4Zqb
jCtFD7HSgGG/0QN6HNpPgWPuqKKmdKgWVBQ5U3+Y7wAQnnqpxQJbBQf9w8Tae30xWhPC+h5hwmhw
wcUQ087irXM/7bA1ACqvx0Wcu+1EgEmyavdemncfra5kprCV/9n3Einbv/eMH0iRs7HAU8EotNj/
EpEBH16TO5nvZ6gVLWSVKvLtsoSkZ8CbeTgFSlNkyCZ/AnyPxWLxsV63CvPbrTUK0sGugl2f+IgZ
vBi2sqMYtix6q/mQNm1t4nvru3Fm2HZ5V1pUJg5Gy//r9kLlbKCByWRFhTdMTe4EAKOeTpRzU/zl
XtPBlI/Pkan3WmTVqUrPQYPyAMf4qsRkX9Dm68hRAvqBGlT8Sa9jJa4Rc5+J5Xn1jCmtJiXEglrr
KE06djtjaJoqlEXLpvvhJVGgEbCMdugzlYRpCtGpdRyeJrsTJCs1IoRyTdMY0ruTJkrsAAAjQ7e+
jZc2T60zQaW0FSb2rOe47HKDgXax1otxLwEpBJy3NLWP4argyTsV3iiWIe3b1eA+T9653UIkDKbL
4q/I3oED6Y6L8PK0TO/CxUEBBekbb9yabRPmR724iqMOEXC03s9SY7YLmR13p98saer4Xu0v+vAF
F6/xjPC98lm5VdJKMGe7xr8zbBv3i8PzrDl0jDQMOpuWoYlxUqLY9STKrKKnn6esHiMVU/T83om4
XYPKPAJPKzJaR4uhXDROc+x8/5StsZS1sfsLgPp6hvYCOOMat7Fq4ayrghwshlFV3qi7D5pugl7g
27leq+mW1VhW3Tgj+6+EVdFX8TavsyRkuykBRz3OXvqdLFcanaPZehvM4M2TG9l34B0UhVIiQGvV
3ssfT9kvL/GCVwW+pP5OwyRMbUnfAqqPT9YOB8V/AMiHgMz5w+LSmdStn5GVBTWhHgksfzojNc92
p7ols1b19F/Xx/VtGP92YVrzQsLo4qQ+vR70gwsBz9eLu5ClouLQXiR0Em+sDVMnfXctoP7CuoQx
i3qBSmnSKOv1P2Hz7C5KX9+rwJuMLkrPIEgTTX8KkgeoXsiBG5gKwGPT3dpAq7hSTuwXMvZ+R3Om
AMrrS5XsFPxzOAsqlDD+sqt51kZd7sQ5UiPx5GqxqzH+W2KT58e/ZpegV57TX+sntpXDWSdou9WN
PaaAgj9mp8dlOTKd/8WLU719uK03NInnbwKlapoalG/VC8pB9w5goKPiLs31HOVmV3qrGFiZZTUX
UH+/O+vci6+xjO485MV68DFzmuTWFPsJ/QWewwbLmQJXFg/13Znhy1CyJ+sq4nx7zmnBpKMY0igi
X41J5XWWYCmeu4LmOGHeu2dVgr7z/EJT40eCmaFSXy/Sncz7GnOcJeh5yN4R42OUsg5igbv04Sdv
y4E0w4LFvxz8+i+zH3JdJZhKDF7l1tLqbdhdPNrHEmgVh5tD5ChzjHx9sviIgLkgdIGwTuLPHquF
iCmLbCQKQk8OnSGC6P9nbRA7kc2KFpdPPsVwDlyDOBNBeJWSzMYiuwSSTLoEAqxCsBx395ItGcWu
lBQ5JJqlUV1e/dnFr2+BI1FZPrFCGNv+uG/CUxvdY48Y0xOfLL2px0Jg9X9AMPKLbmqoljlFLYZ6
jX5EhWaLXAd3kpG3HvCU6EePtZQ5TzTP9AqUrcNpXEqGAyu/b8uXbzMKcZgKRf2Wfb6bNqf69v9t
t6wAdXZYF5zlJXCyv++cdbKclSda9x8MF24l8b1MQwlbKC5cZEaqdr4TA9SStV07bdLNQDNphqCO
UvVhbmk/tC7w7iGVYhZx4l3jZEUBOGDxvLXIATJ/pPYDmAczAySyHKoSnsT+Oi+lhpE/rwwTmVcQ
HkRp1l0fXiK9Dgl/klVkqMN6fI9habCnPbLfBqlDv2YK047MbS/Zwzxo1HITchWDtfYalOJaxWYw
ogXC97UqnAY/i3Ub7MMX0I0avVx1OO88BWZYWIfIsgJpJ4/Iy/2LdjukL3GVI9q279qT2jdwBBAo
Ag6euzyCXDkpaLV9qI5kXdUBU8jKoyiwSS9IRL1XAE9BNvkh4qrODAR3cpimbu0nZTgxCPu1pT8p
KhVesisCK6IDtzJzZ2q+O3LtNTqpnYFEbuTw01GytwkEWRv7k3YxMDJXXT5TIhTS0/ADsrH2Fw1X
y83A/qlkwRZEDsYs5W4Z9YA6eQJ6WeVwUCuxNy9PQ718gL7oS9ngmLoJsVx180lgvE8r6df8MFkp
vimCS+dl/lkn/IM/5buQ7pSbzxPXA8tWXVU3os5ejpgCEXh4GLpAzxQNpL/+oE91pT2okCXDVizi
59asqqZw7DU/pmS142pp0N84vdPd9MDqEIlhHXw5054CVfTYNkr5GHqn6sQ8Ej6aa91hpjRI8zF1
0OIt51tCYyzPd0a4jnNy3uRSiOLZuPhofOvjLJGo4e/oCvTL9w1tSYlY/phYBkwRWeAUshlfjpqD
DMnwMiV7jjDryinXWHb8mLA0kwFX5sPzoS4evi/9Sdf1KbBASDrAmZYFOb6AkY47uptg4YcHikf3
sZf+wXDLNi/1BapVXWdYqd/aNpkZoKrw0SqY84ZGw/dtoGq9u6EgEG5FbMH7EtZbxh1UGGpenVev
uPKY+fhHZbnkryZ5IXbKov6fLvxTcZ8UqCHEzMhDKFmJfSoWJYpFvuAH2tMN7B1CKG6Jr1Ryb9PI
Av88pD6amXo5N7z8Jc7FylREQWa9aqiG7dcOb5XiN0GLeJJa18vEo+1XOsfEoSYM5fbdddXvDjSs
Ft67breYKMPfMuk+HZlEO6N5om8SEH1LbfkoMhRp////8I6lqN7RdO66jmFrEKlqOo2gGpbJn3h1
BKnPtPxvwKIbrJVU6L17H1aEh8NhKiHfJiKIB0T59/39LEyEbZJ5oENYYAbzqqOjuWuwsLZnrz31
d1IUjSjVX3gFZXdloHhxorKSz+YKQqmlgTY/g8Uco8+e1/coJHN/GFmbeUkf2sqDXnT2ZFn0Jn29
mx/mFU2WpRXbg6P8g3nFYyqiPJgYHZbm7pu0qFh9nsznN0KveJvigGaeSZd8EFwWcSDMBhO9l3+F
7FE3kectJ1h8o8rwT/l6Bc4BWPykD64QNE3m0mVPTwsDbOrLS4W2jogM8C4o4eUN4OiL1YxNUprF
UtzVKAGf0iwB6awBNoQtAZTbTGTRIKdgBfPFCbot3lbtaSdpN1UrdlNUFvmn/mN1Q9xAsO4Z5fA6
v+90Ht3jJM/A01h09BZykWnWRYTb8Q0q8Zq8KfXh8+AebNSILw2B50l/VeD9L8bVaiqPqL3rF6BG
ndBJwS9CFjU5Bmp3meSeb445bVBPjeXcwiqiQVO5kIf5Fj3ZXyf+vTUKMM1O7cttFqjBB80QDZ+U
nH4kgDLUsmXqu5S+65ZOCdoMpT9Cgm1iR24m2BpscNHUKO8NNXgcYTg7aifOKdkQUuHNZD7CwgMz
Bie87ddxAPVDU9u9FFTi6WgG8VPj2ibUYr9Ox2sVmNDZz5o/YLiNxHPvdQ+/jWd/XDA2tVvyltAU
iHlaw6CTi1DBAmmb6qGUrmM0lokQL7arQdDx+16OKRgsYutUlPcHFCAXSJOXXurhTTNTNDMBu4Sk
kGzh4x3/lDZzK/cqg47SOVV5HIZuJ+nRPqoW+fP8tiob1k/MjXn7W1hCH5YAxI8O54PeSeDc9hXz
NWIzRSrQdrwH0mqHjQ50uJNAKdH0ls8Gz/uu72ridr6LSwW87ujO7lpcZ0T9i4JM9nzBhzWuO38M
a8duWugb//4HAKD/Fll5GRJVFItfr8069aEYC2d9zth/8yw73utXrbYb4eiZV+ltVfYnnv75ivRB
MQW/D6jwcsDsBR9f99PMYjM7VCHq0P4WblRx0vY3ETo+ngWFR/Zor8cTnkV6fcKylG6Ft8ii62In
/3FO+RlEktAIzaK8muOyx6fxLttb8rwFA/l4N1FN9UrvqhHmj7Ae9hjftgnNy/n0Xf/tmSETc9oD
SIu5lbZWWY3oGCf6llZxhwZijChHJK5wMhC1ck5gA/0u6UyVthSLw+ges9Ko1/MTNUFBHQbpogaV
TT0ZYk17qgPeavEAf21l6KBOLf+KcYA7phSzTXeYsZcVIADo7/cziiUwWlsVno6I3TfuQA38R+2i
MT3rLuXv/32TkgNFIGwK3vP1UxXV1jo+Iw7mUsiZVk5jK6oUMDKqKKS8LKSnBJsaeUXOP+AHyjRG
cVlSD1mJzst5Ykc96bZZXZylBf/tVXuE8Mq+6e2XOA/0HlyrzUfprECA9M0gOhSP2RNdFwBRhhOB
dmt+fuCIyeuxUmW59IhJa0Y5TTgFyG/0eyFpR2drKRMzAIvWu2BDTZRVLJvtzGrwxOzvLDzROg65
VTsYOen7AXvPJJgkHqiPebVrGApKM+dqUJLg2Wt1gTE4XXOQZIcF0eVBLsC7y72WRJrtEufSfrBp
qfWGkkqG54F22pCES/dimZPC6YxgtBslNJhZTgdvIsZRtD9xUS7hRJRxqWwfQtBYecXhabHESWac
WYrgC6pRExyIfgGpsP+q+J/V7KiDGDeff7/0zFyWDO6rM8rzmyQiT/25ZDO2xoXfqkp5SQGnhXWa
qZyhHx8hqn8JT1whevsT5WoWuOteoElZwjHnAXpOW/OxkeJfyVVS2I0WaOpR+Ep5JQeYPfDOYMJW
qldDP3z+f0tK15WAQcthJGv2jaiT5+xPX+o73Jm0i0Kcmnj4rxD7fqWKirDgtTAL1elyo7gmesXQ
3QR/cyTgcIFTkNAxwuN+4ikOcL2WmLdaTDuZWg3lx8GCySzF8uwZmPsFsF9odHqeDJIY6aOJ0bF0
YyYnjgY4HVwx3diOFtnfiJlEQTYRP1UfOPIAo8LMJG61bZmN9pIeWRyac9mPN/q6RLk5/NBgGW9t
EvHcXQk+eDJZXj0qnwsR6Con7T6U3WVgsLHsbg5tb2+dfUfu5VfOLfstqkAcE9x9keFShstMX5ps
gL5OcjfaoGjBooBzD8O31tvU66WvEKSJq2UN4pAN7QPhr6VvEcNv0TZBomhqnO+j7tz4Ai1+ZPaU
ff0UVaDnYt/5LtkBXZgxVJ1uqY15SwBxfVEdqGSlgX1EZ4Yn1RYTbc7hmxM/BVhzKyPWJunr5Zg/
4tHR2duye1AgWJz8nJgmv4EPQTU4b0V0O1s/5Zns9Gq2r82EDF1Mt/BV4hglG+UYdUlw0+oJKaw8
cq4Y5FNBofMnOmqigX0RPOag20ZAg649tCXuwgWlk+XvyBWgIAAf4nYVbMr3oBn9TNrx1aIrHfap
QJKVFGtkpIEVvwLUHmaEPYUwP9pAk75D+KprZeEs1dT+s46AoOYKlzfKyOZOtCMush4wzhYEh/nJ
mi58D4Lt5L2dH82FNxdvcgltUkSN5cI2KpE3EMy2g/WkV3JprG0NiW9gCAdpOzYoSoH2+RxbmrD4
GTEIcFrwtxteI/2HvM85M1f8HRbQ4+7LjEiGg+g5iUy/wdC6jF0QqVA340zJXHovDmjhvOMdIxfq
etdg9QrYe7YxtIE8+DsenSD9vJFlbPw8zF4JpNtGvfFHbj20acTdFVbkT/r2kVzgvEJdCjdllney
3CHPLU9YlWyfIz9i2CXAzTKE7tm9zPifHiKxTYVwz0qqBw5GQSnpAyD57pOj0Yh0QekbDmqa4t+8
9w/GCn5RYMfphBimkYWNsE/h82i/Q+X3CdoelMInXYNhsgklOYoRwFUbQEDkI7Thd6H6VMXE3I3K
yP9Ttue9CGy3Mm8CZxkpkqlOi0uq3ZpA2RO7hMmkzqa6IfIMmkd15iGBUexXrNXNdUb84pVGhD9S
NixJKdb31TTtrcS4YstlgklLzm52m0bxY56u5vVpsJ2wJJQ9G9gPje4D80eI4LTgKFSuxUtuMQt6
eb+Y7+bLoiu08GP0uhQLz+1Ll7SR/l2pFeyS/1eDieiDW12WUVXQzKBcBrNSiIPttSSO2mIHL8UK
uE3sacmlksXoOPGjmZ5KZvBkqS3epl2lZCmdO/n0ZLgTAhwKHtIuxA+e39hO3p+tQnXTdfcfchIv
kG2znH1R+AjgwWgj0K9UEl2uh3uf4igeFAfq+4pFg4rfSMOMXdbh0+uPIdQCUbUcgAuUjZtU+nK9
34wF4QrTqoYtDarHBZqGFFz7jf69O92QvgyKXGkpuDuAM592RfNLj3z2ieecv2YDezeZP5txxrxh
KF7TMANsGVyGG2enV833tsf2o1Cz+WCqw61d+vWS8SUKgsxrO+GV+3t4+uCc+P5dAYyo5aT5OCT0
yTLapYbpPiuEHEn/IuwnM6XYuhWYqTexLBeBWU4hk3YOmtv6fz9xNOoEp1cTAlvrhr0tSensUeq9
O4xzGCNVpoybSLG5Dy+OLJy87bICOm96NTyoOs+pDPKzVZg5ol2wSDCOadKzdmD9DbkbhTgAByUk
69qIfBnuFWNLJgMH4zcgg2Ak19JLKHV2fylLcWQ53ASyZpaDpwbxTl7KTe3YxrWBO43J1RbSt3jt
tX3NXpkDnX7GDKWp9cUoIeBGJMuvUQ6SkomTST01FipRS18yGcy71FSAhNB0Wo+z6ywuBMXVNK9R
cioVY71WSPZZAwMYHYRp0L4+4UOvM5u1O6yZZhJRB9NiOCfbBFz2CzaXw+oZHahQqJFTgUwpGqpV
lI8HmeNLo2JmLmu4DEy5iRyS4SdrxJ1DFHg1b+xVeAaZphzCAEj5uOI3PTmY7N9gvZUy0KP/xJ1P
KzORr4nksLGnuIWUeE7TlDcmNon1QP3ubl356kfHPM9HrcCFEK9u2+Qd0NiJzFUB4v4001wEQlN9
aooWST2VD98QT1brAe7vgwbPcOiJk8R3pnryjuzueL8PiSXgFdPVodLa6mJeYtWOzwBgWYRxpspw
3uVWNdzvtEHF81MpWP0E7b3utFwGhwFbre3jNUGvZwwbTEeqYZFuLNGZXa4LS6zMYAPSJ6KfVPTD
hQXFYXelLhDcXG3x5BQlAhPdWiRPfQ2NefW8zD4XUT+7feN7yTKdM8RCm8Li5LzJ+YB6HDkIIlvc
crZKjsLfyLcHNoGya2Z3xyhuPT25k7sgXOz4Ht542niv3H0DmijAjcMTTbQthIZ5CT+NdAPFaRQU
TyeIzGaH4k+YjhFXNxyCREEBaQTm7q4pxBRYNSseF9KVuCT1efwoOEYI8Bdwz252IfEJqTGB6MXz
BcZAcup/m8L7rIcEtjyjCfzmiXR0J7IFQvTgkL1qwIw7mmJAqtXrYxGdO+BRVRMZ5zqATCtUPNWe
CBqoZv+qLquzU9hHvPVzpq98/vyiyDx0IkYAHVvJqSv2vXTM/cnnBma//SWQDHpbtHVjImfTa8Sk
EYOe7LAKJBCtv7lTq88A/U61nrXq8P4vcJB0knH2J6FRhQMw/68MjGv92UWHL+pVobtvonoUGfNt
EbuRxfi2sxgQDF8Fk8DeC0JPXSomln1CsFSqfSauQ3rK4n2bHjeaAb7R4ezcx3PLrg0zbrho8M73
1m4RPAHxwzKmlozi78a1Se8qJCVro69x5dLBGOKixxW0fPPz084/OQzdKep8fShs+sLuKur4hu6K
VsTzQhd9VyKHBzZfhzUgTi4cPS86jEoYB+LVlqrU+ABDCkcAnlEiRGC3PAtGu0wwZ12jnBj03f4R
1e0k/qhqIA2t5CZDNeAoK3uSKbFuUP/ixjC0W2tmS6WPJfU//tZ3gQbQByYm9+24BbE+F9Ox1O32
2TWapjIT1Bofa1ZTQyWFyyhYrhzcN9xX3qx/f5RYDIyhvQkH6ZWbu+MQxIGC17GMYKcbpe15He1k
zrK/I2174ZsvjXimOIrwY0NLajaTsrg5gEZHQ4THORiqU+iZ6DPGRstDuPAmxJpjU6RIi7L8b9dN
SX0k7YtpyC0ZYwEv8c4oFZX1OaB54pGmpfYGrTwreQPJl6u5mwH/FYqFfqKXy03plo5KNMnWoZS+
BDJZBBVAWtuEPxSga/6s/utVtizWTNE97B37rdIQhvjehtazyL3YUXcKS77Xy2S7K4ERwxKIv7FB
6GWgY4Dcjtpd8aa7mMIfYgbi8VlWPaA5NJT2BXI8PGLkqLc4GFxAhY9fpKAqkxbpbczjh06k8okD
WCNT5PvacugGuftvmA2cGOeIwKEtz9dIyoRijRf3RuxPxESvg16EAZ2NB+Y86myMevjB7VR7KIKe
+kzAI/ln2iLw/F7YMC5eQLAW9EDYzeXChlhdlX1SI9obJTXeO+ztS84sEDEDMm4PmJx2RHFqo9Lo
sOM07Hfv151L/mutq4gQ2RKVV9ZME4CHSKIw0++wF03M4+Z+3OJvB5EUwxkvRjKv7kcCsf7Ol5LL
nBJfqTGtKglmrNwkp6kKFymWnTiq2EDMPpsVSZw/sypWXACq+JGWaHhfT2R0AdZk8LK2/qxAFFGL
Bo9XqbMghWlF3debnCudsk8/2i27fKbFt6pYGWVQgKYe3lIEkLbdohHkVQuVBDaWBx76ZAYU3tJj
IA0AYT7ybginNjOfGkpXE+BpUKF3rjhg/TKKb6nbC58oTw5tMJ4iUpmgPRAEpkPeaGtW+aLDbrUy
bSd4UXdJTInjiYTlAMWxF42tIm7mtM4hr0+2f0DjFNeOtemfhCI0I24aKXwAUZonm9R2wAQm7k0z
82RndUUXZU6HZNXPopvu1SRlqYkmvI0gw6Hblf6BsZL2pmVc5mYk62836cbF/VvteLAR7XfkwGt2
pdkDPo4gbRThrGZVOnMQCae98zpW4UIEBqbJWmNlcCLDNcleo2qI9rsuRhRRpEhiwGdRG4IEBQ4B
B0ljTo2n0azIQe0sfEEZY05boIqSs3gbis8k7TF8uKCYp2XreATa7Lra7RcGdBFk5WBUa6jnJu7t
cYjkI6hifa8+S2WQgomjipw1AhKtW9/LWMAwO9hGQG4kQ3+6EQQZWI98Cg0Kp0iWazs57/FbPVbr
5l/VD1cpvu1Sw3LsM5hC12ioOEwYQHxb6dXgTmq60RA55IlN1wvWYfWNeTSlf2YdmsIn/VtYzRDx
1eli0qNa76w2sVuMvcOg0XsgIe32IHpy4l8PfRAmb3jbbZxCB8kLUkQEVKt5SazVOSX/jmYP/9+4
xhjVDZQZVL1/FIscmoL2NDPfia4YiwF25LzVvf755dmETGHVDhyQtHwJjewMDyWtgV/9FaSRWJTW
ZNmCq6hJwGO1gYp8hN/wibCPL/xG8WpB8xP79u5+WCYR7EJUDUnTaKB5PYwZtPnX5MJne8zKqfH0
Z57RMPfDmUadphOGutZcs7P7p2xHNAQnpF6Rgo+8aiV2S/sLUeSDWBB3wNYA+eGqBRyr+kKuqZwI
7YEj6SXhhY93IgOgFhmVB0bcmYpxRzCE3LnxFee3quL2mVcb2QMYq5SIQGQnGPQrVs1aigtYt8ep
AKMviXwf09M3RCY3bLhk57A3UTiQgr/XR1xo293Q9KwoIMEPzWEHwx6najGnlqgYHgb3Htf/QeuW
R/wpSG/Ifjr3GpIxnLm4W2UJNtrhfzXcYkc/trCzrfzssPlQnx7frgTYaEap3FGj2/t6wVwk005z
RESnKoUmOjmTenOn2rGAeAuC5bxt1/caPtSDOYSseXQVu4rxV2I0CyYwpgOxHK0P40J6I2b8tlcv
YrulhevjV1PtF/q4+ZExiZlnG1Mu2BAr2lx+keE1nn5On85oSQiHlH8ABASHVZYxncLW+Kkvnrr/
O6A3hI/3oEPOBmCQK6ta2lTM9OmekJDHJTXXTvEJ9j3Yd75GT2AZhvQoy0hvFzWutSX1vEb3OAm0
HIxMg1fy2uc74d385KcVCPekb6sgSejm3gg4d/woLMSgbme3MyJqflZIjZa35vuT9Lnm5gJAlbtx
XgXVJNBdX07n5KLxNMJGSsSAvSfDNIFTAuGSZbYxdO+0Hljnrgyw1ogSRE08SorewlKJ1tYFUaRG
Q10HNxMJCoarl2AKifQDMLDaa2Fcr4gsObdTC5echM4GVQGumYCV9amrjUzQ+2os7p67pH6BPMTz
/qobYvq9IYby2WxNH5Eh5yU+phqdU9pxcK/xD03BDZ2liarBnNMt3Bw5c5Pnt9Bx9MityjTOclnR
6Y6j03M4jUXazLDLsRqlC7vl2ZFXHyX6HJmeZKxMyxu0u5/YngZsx11Cpe+wfMNoR/3OcxNcW95M
kjene9ZkGpgwaS1csNZD+cOc8VJQm0sNtnHkNEFyumr2bwjB9A6Jf2gd0j7qfFXtWpvDz6J/N00T
eizNcW+qIToZQOYOogwBqasFgdm3dNm0iYmB3PznfjOWwm1GhfqrlPp7nvl9leUx82QpJ7i0lNKm
fV9kQJ5fYdmLAc6B+UoFVBjRS3LumUx0f49wfN3MyL0liI51KSEjU4S0Rv1uTTKbNOric1zABW1P
pLCH1GoYEjySoEUbvj42mO77VpwkFK/z+u1OT2mBa/tpZJKdbhRd2roDFiqM+CRnUrvB0431r1co
Ug9pA8qqkDFsbOLZEPzbiQ+7zzC8VHHLynvj3rLz0wKtp+ntjJvogxEC04wmEBqC4CKdDX+Bl9n8
SiPlYNqVsmrDkNBONhgRDMY3B0/Szx/erobrVcff2AaIIyLM49z75tzfz7Vjja1rRa34EQLaCcSd
q/GGBG+wVjIY/eK+vNbQFMXAsB9f3fhAPPB9W6oT8s08KUm59EpLzBXZhrC9v12l6dtonr+c0+DM
pK2jVrHo70Dac2g7Z69udtaQniUayUNV/XeTP1GxV7V7xCLj355lmsAUQUzNmo/ssO0hYq/pxvxV
z0yRhUEopVWaVJmN4g7yCCsOtGKybs5guaYEK7LxFUoEpNhtiwPS7xl5jGHeGioxXCMtRNxL3MIK
Ss4+sfGtzySw5pzZFctj9F5aAX/X93uMHOrJM3YgAUb4u6oZJ2uXrQZn0AdHqwvKNSiioYIkF+//
SPb4xsJn4Yr3z8G2eykuqcUg9elWXIxev3txml05o28RpyKHmmj//DLoXlkHicbK1Y4mZTnpDBRq
lHWyqNmaqHExQ8FR5PITvs2cs2Tg6BHtXVYHukp69Pfn81bzkgNQTB3ObPmQHUsM0V4IwwXyieIF
GK8FNQr+QcaTHVVQqFRohGNm5XVBE3Kc/axv10xaOwQWd6ygqbWVstg4x5kJQZRe/iWPvogUiXZ+
kDjhqnz3xV2uczuge85gjrCh/7J2RpJ6hIreXpkrn9Eb4fWXjGJrX1/uZIEdpRMXzW1ud9XIobq8
0YRUCvp5ix6a8Wt7wlCMqIxRGozR758dc43o6X9MBnrrUlXZlmXTGnvjtRAg+VGTx3mwmKEHNEsZ
26NEEv4AFyU+rttudWMPKxcZErSpkc9KAa0z40a82dukjntMp948ujzij0pGfD0a9jtXWc/d/rdA
MHZnJEs09oPCGwY/wkF1IEjhAG2gpWGkOmqgsUwWXhLyMBHK81KmAo6sPiuDK4vCKgD0vATpvM0k
RTG2AkAv+wi4rpILK9deUJLGV08e8xZPEV3FHC/Ys3GcvMsaltyKtnDISv47EpeSiPTosOzjvFWZ
xK2CdKetnGTGOunNgASeVnG9Llcg5JSineu2kf/awmNCJJFdahvFspMoQNa9dOOW/scTHqyLyvcJ
o5u6RcxO9z6OKTo7DeKB6ve9ofoq/JUC/yEfkuTtHfg3ehWhoibvfDN7KAp/4taH0iQJfxMOLo2Z
2BKrVMnASM9J304/H7po44FBmdIKxyC4D6BlCHLKJgtHghbVS+LoABZ6qqqwPRHGLFidQFOFeeE6
5ketS+WNdpX18PX1R+4MJr4tUjqTM/FVy9pNbxFmwycIfsXUfGOMiOptN4VXttjDeopTk/Omjwye
R7ZWiVn19ssrVmxYadF+0U/6u9CGoWs9FR8Sn5gDwOeVuyDNspqTcmv1oyfkgefGCtAWtBQy4bmU
PZpAr731iB9vWONzF6HvTi+VhQaWtBNVkZDjNRv1wPTx7IlP5+RhJgqVBXP3lBLacLGuZtCZ4+ko
raZ2qUY5CE430lqgEPNkLP5oQSBsxnhKgsaL/nxMYXRHgw0OC6Q+FqUmT2PX12LQze6qGGIZ1wFQ
npzcGITQwpaf1Zz8d9LfOj199ytkB257UDE4p+nZbRRKWapJqXGiyAtbwyiTF55E2baWClF7mnHf
D6voJLyzpNaP0Jdhc4Bj4DsQZtZZUYg3z5tW09AZd75UIREwtAS0WoA2NdqVo3zjjTn0Ss3yt5z9
DhSMr6F1YVgwO08s4EOjgymZrFVHd5/MrYf0kTfOFXYgXUNDMA0d9LZWPdTRfns7bcgdNMISLhHB
tk7TgYI7PQwk3H4CiL+FA9wG7CJjv4CBVLqMxYDcD5fTVqQvmkA/1TV+ly5W7Ck2WpuMpDjNfaq2
aUdDgYAI4W/Fg//ugJc4lueCJEv250dUIpZkeVfkC30Eh7LBx5EnX66mEfqOPRKUBe30N1OZdpW4
+IJ6Bj8bMsylxl4DB5juIGbXSJdELtLHhnnE4Rd0tBvLoy1cTOr1Vif3QLvjNCbo9jiXgm9J7MOJ
T/ONaS04aS0D0Q1nGEBfnc7Ucd1R2zdXhNdFQf/F8hHp6Bw+9yWzPGL0R3niJUSb2+LC5RHxnLq2
pwDaaTSXSAeA0cSCkmwHvFH05fT9CF+uGr1FLM2emfqXN8qX16X208/9DnHp4Vu9RgPTsa95Pr6e
4rVwmTRaUoIDtzyJu3dcKlNEaypj9P6rBNFYBD9n2T2RAwiYnsyqXaU0LFx1uiu0o0umyrhGjLOr
pFo+WyhA0XtRSSAZmVXGjGK07Mjt6YqdKiarozYRM0NFRf7O6V7hh+i8UMoE/BV1SLsL0lHNRYr6
XRwiJNqPQzUs3QqapCqUuSh9ipy4fU1YuI8Ua3uv+cmDgg9VjoARGMxfqFlsPUM4D1d4tDRRDWC5
GwnzGS8PV/ZdK6ik6xkbRHqsDefWzS9hMUOruCNLjVlQuhIm8RMI/Y8zwhq/8VkNvpK8EgppPYcP
g2wM8Hl+WKlmx22Vo7vujjNP70u6eBsAK/Vv+xvow9jMvt+T7FCAQOHn2N1WPYfttGFvydmAsK6S
hSQpvzj5kqegNEOOjbCiBhaga/WaLsw0CINxGn4Q6XMQN+Gcm/Qt3S48Tg/oot6eRJfgxcBMAb6t
AqHx2ILhuf33gEItHImuP+e/PmXlT8pCLhoortQ017Chd+C2CTXVLZngOz3TnE9MSknvWiEWO1jw
uPXmt1W/zAfiAbxqafEoLa0qP39rFP54xFLoyUTKWCZ8pAxno7oI9KonMEnHfYfbQUQmmSL9bumP
sEN9a52F7Id/9k+apvO01DZrvARKGGsv9dEqEQsrGq9nxYnzOc30K7xR4ZaZr1xaz3CQ9E/V0G+U
LMx9m3x4kAFzyRrgUyI2GgwPIq67L7+jnvaTEXsXCeWnTISPeW9LGzicfKJdaIns9I7oQgahTRGf
sclFVRfR0riQqJi1VuUu6FeptFMX096vuIfos+6oeQ2MWP5QoAU4gOcU+zGlOTJVZphWu1FMpLez
Pju3S6zmbRTFVaFyvxXsV3IJKO8tNRTdRbH5nEVo3xaZmgx4UyaFgyk9lwN1OLmtxmFcxLvQk/3s
+SibbzP37kXqZEfpYFgN0zmwPnS2qk1u/BZ29pYGjoQGFdIXSQvYSHRaTMq/2Uj4UZcBavOzQ6r4
BC0EeFr/oI3jTu2nRP7BsiMIyDXhk4285WYHgpkZOjS+ULL7ClOMxO8zBkwLNXixZHTZAX+c2Sep
YyLovjUoCzgXlArFtvL+b0zaLwe6uv6d+bN7dk+e1ywF+ZPHkkYDKmUAG9HMo9854/v7bFNq1KLy
MqmhFCJqTzxxshy4NwF2kCCvY2Q+H4FxXVy8M0Z1YbWpKZSp8djS0ox8FhS1bUyK4eMdmvVjVQS8
P2cGvpIrjCFP1VILvLyOCTLue8UNB4t5IdU3DEWJdt9fGS5ESP1/Uqj3vUhM1KHaOaDjxtJpf1zF
z8YmVf/+W4wt5i4wldYaloeo3+rgfQSQeErC60xjHu3LKKFlf4Blx0janxluWUAgX0gb4AvseXn2
kCBHhXJSmcyIjy+by+kCCBZE1EDagXSGKHyDYuDFlcc/kzGKmb/FsAd8Z6HDYkk0pSWz+0eseNih
rNyl+c05o7xzejlowqSmhEu/GYWeC3Sbium2lY6nOCDUsLN4S5smvRybxcKFLmK7yyqL+YIbUBfW
Z+OllosYwUWFvcjWiUd+NXNZ9uWeI0cFuvA1c1f0i4wmHtU8+nypRgrH2OlQadHD2uOXzYmdCz1q
KGKXJRymfi299Dyn9K6xtMiL3WcAK1HLp+RX4QxouRT6W0WAPCikn1JkHAS1V465/C0H1i2lIdPV
A2K8A2XAWJseajTmPQDXgFJO1sdEyMds8tF0Lo945/Gffc/xai1jzUv8bm0uAl/ncJaNKZugdtwp
rLd4xEiEogcBJguZ63obGyXe3R5Un7513p7s8JMzAd62XtIb8oFOF/QjNkDF8pux1RL/svbpvsga
KfGFOJLjh14sG7PzEVEfMgF1APexwY54beQn4QjucNNocgFlLTMEvWMLSI2zaYyjBCBZ4n6zv9Vx
of5TR8ZhSUy8Lku/Fw7f3dGOLsHG9r/g8VUzzCIKou0ZE0wcZqs/Lkk3XYVkURKBt5OWS1ZXeU6Q
MQDBVqK76yIBy02Tx6U2lysnpS55Oi9tkub2rjMOSYpvlGJjUKlc63qMyr2S5Wa52y5GyJAh068G
3T7pM9XGW4iHd+dqQoLEmPgb9+WerQNYMW4sEKZEAyPi6x51hy+0k8ogOp2q/Wz/atclueEpfKzE
gaMsDpHJkXrd5rjpi9j6rWApasCLRKKjmHQqqRnrCT8t9gRhlAcdKOkniHBcsTWtDeEHT6hG+Jig
HPW1N1bWIle3bOJOfMcEHrfs6tX40P2wl5XP8+heY+pBEEeeQs8OSa7W8Nbw8SYWUPg/3CbBI8Dx
aZ49DaAU9PfcIYNzPcpTY3cs4CyNw7lhZRHRC3HXLcJqZQiO41NmhTGnsaJT/+5+GsIPrROb1e2J
W1GNh6qDMAE5qkJyjc2kTceyFPQ8liV+xrPIPhZBqJ+W7wju+8tYr2usDgIibUh8yMN2rFrGVFAV
3ndobpRgvLJ6/Upru4nUHEL+0hP5LsXpnOCanUhc6hpJVxHn73W+AMrnyisN0rN/ifVKBz0l+Y/9
ltJJVBa1UtR/BtAXVpudUDPAumXrTGAF5ecX7NKIcGeU2Jz0h65UmyRhoewKHqNfp4oRttpll2Xk
1HE5TKQwE20nAMhd8kdbUXQsvojRHsEcvheIHOQ6wRt67EBvLxVic3Sg5IlG2grAR0/1LZ++6BFD
5+2gWYcw662R3wcBD8u1sN9Dm0HEKB8DMRPgdp/EqdxdjwffM2bFvYznBSRiwKkL1us0ePOQ0IK6
khzdasro2FDeLzG08kL+BYTOv9aDYgueOObEbq1e8PUZsUqiYQQkp4lKPzQKYdWlMlWyOjoM3m1G
zoDrFYiFntLX+RFrhnR1W1OHPW6Z8qphbvIHeMh/e9/cOgDzpEotVr4qssMEIe1CKZhm2h+n0kUn
G1Q92pOEQYo6XpMLcgdX3C+WXuwzAjZBj3NFc7vG6HJ0s1vSLcC1BBtNnXXTsfefsiz6O21ZqBo6
CHjjsLE3ptmp/tI6BWadmlkxiCdCuONYnqORuvv7K9yWGLpdb9+l25xapqx6ag8hR/CpguPn111a
A8184wZErdeHIM+TkKMJEQTssPo+BLSzKdF2xwM+MlwxnIPt6yyTTOQzVWC6r/7G9+EhYPNQ6xJi
XFyi2AW9NzEoiDT0cmfBrgAG6+Xko8NjVxWwRuhyZc1IjsHs2hb++R8SaMK41TLfNGKNO+S/4/jX
aQ8QH+wcqwNGTFP7bXKxTjA2BokHiH6Or/fg2bz/eJTY5z1leUJvPpk8uV4iBM5M3XU53mFZt+2r
43hqO03NqfXfxMsPQvGsRrgByDyht96nypdo/bvuaZwkwzxl+YVm76rhRE8gavripgpSjuM2C8/Q
QG5yOqHvPkS4YZQwzg8P5wQhSk1vCuAz9AYAsWht32oYae2eJfwoioNLpDPoT6HNyxjM7xMttWhY
7RwClXuGk/P8dX16Ucf8L4J3XiUtMqQso1chroJq5SlpP+PC9R1Z+LCK4H2JMyDQ3p0th3Itaw0X
hhs7bT9Ag+tkKhBca0zJ4OJxg0AS2+0dMuRf5F/zek6dzyBdu7E/sYjlLNpd8mbgIDK8VMgKv6kK
VUNDQ+oBgcrc3wSn/k2gn0s5hyc/N9XE8j7VEaV2UkQP/MwC7ph6KQLskw0f+eVnWOYkP62K3tif
+mrYno0nG0YpoR3zoh0wlOKAhs9nCZmR9+XUNrmCEgMa8qFdlcc+5YaRKxEO+1crNUaS/sUgkiPc
XZcoVi1+UU7dCHsKbkIFTrVCOYsqckPJeFVbGODw6hMtOkyC5PTdsNrD2fP9x1wG9OgCUvkjrUYg
+QADXncRcIgfoIkEdjnMeiW+fRm+MG1j0NwNaAuOOoKEBbVCLWmAPCLd9Neri38+QX+Ll76WHndp
NeMA0CnpQazm+tk3BnoJRa6pcY/gQaL/vDm5pncnQz9CrOOVxoV3hbrr4C5OBKIz8/dH/LegCc7y
MUKevmMOw973MeYe/z/MEcUtid+KNn27duKXiwIBZXAlbH2maY70v+aF8MxEBMJsov6kDzWjU3Gt
fnLcGImZgu2o4lGfMUzFRPDvoiirl5xnIaL3p27e6mJPpCCdAtJK88PAyNBr9l4CP5Eo2i3xhaeP
flLO+YnkOReMjCPyoFWlpFwlD03aN5MMYchjTVT9K/knHwSrTzvE7Q2QS6bmvFgnRusTuwdebLjq
6gb99g2ycerEFtV5onLfAzsQIkcbRJAE5hnXrpjyMBoYcz1fT9VhO+f2iYGiNFQb5DpL0y3Cy2ro
V1/UosmlBhpmIjk4U/cdXiH8S3pJfkMausPCh4geiJP2koVcmgVqp3TPn5rLjjhZsNzYs6CIp4xL
Cx6qGjII4PSGpXm1Z3jMoGySEajeEAAT4sTyJ6IMjteInWJyGOV4ptRXjn/alaU9i1/BPaEjtiJZ
4C1SeMx/aHZyBhM9lLR9iXkpHRT1r3MpQYUkYKBtXSp6QZ/eoBtXcnDnS2E90X7k0y2D5exAoTW4
E+up/vbl7MDKPiP9AMupA8f66uVfWhqc3rlpcyf8HlMu8ZOWG0Ilw10QdWw8km+22lascygfaQLn
pzrGU4Nyg9l3MdXKh90AOPedqAZh9ZWV+/TYwqU25CzlNXbvPj0IwxjxqlS+uTq3GkrONxjAJqu0
IAbsxjcDbegToQ+h6H+6rgd/hOMHTgTfcD/a+84RP/nd/HuJFZGK7qhveb5otzNfsFs15ofnAPp3
F+Rsw7E4/Y45W/QFdeDa4ZTb4219JoWUMpqZrVWNS+hlrcA5C20xiuk8vjKR3uc99l2BN7BQeC+t
qsPXJwNGg5wCt44bzvoUBuZSBlem3gndBqntK4h/pDYcXvewjjBkA2CpbApaiwbgCJrYVz2kuGkB
Alw+T2+EMoPp0F6SQsLZY2TNcaz3JDZ4fJMa92OV0jvBHOf+Tb3P4gD1oZ2he2sqoOkIrZBwYUgb
Sw/AABIdr2MCtliwAQ6MrldYbwNl63BjJz5Ftb4PE3EkAuhpaSHaj/7zzK+vQDk7vSH2G/t7QzhM
fPhYA/WAdfhJlU+gB6XyguK1fQvtRGajadJZEO8nYBvF++GF9vei0l2E76Q7dB0KjWeF7y/GPewQ
G3uVl8HlXtDAZW6BzoSui4Ytm7LWzlADJhhxm5iD8lbad7LYEdqvPqr29dEZJ6vK4pmmqp8o1xz9
uGolONiJokTGtdk7S8PfhmEBNmGhQUGQyz4SeWDjxtTLms6vaGTAOakTVpHm+3Mmyp+cdof+jZU4
3AYv/7dBzbnTzXh3ZJrCTq1UVhQr3aJiI9UyM4w+zcypFy24vQJSYtlFFlnTWIaknbC5GrA6vV9S
MZE6RELB8zjdgBc9VVoJA0IYGSUiOzQNhEyYW+fXoekulCyO4w0YmFd9KDC8RNLe8W609Auv9YeJ
k8IbyxvzqGVUXqMsZ3StrrHMKPh/Ej5tGJMI1LXmmm/FGf+ZTiII/xuvR+TcvJj3tr+bEW3B/pvn
E5zdva+W+XFMH4Z57pOAGUe6Frgq3T7m3roTfePNQ5JaX7xdZaU65TTngYZ8P7jKMGstwIvt/piU
XKGx0lnRrqABhugolShVLLtky/n81nZuPqwswUuka6p0MQYrfJT2lAXJg6b/jgM/eBBDecUrWszP
xG71nOT0twt6sTxrAzQ8xXi4KNIde0WvF2JVvtW0ykScxZo1kyjsrGCDHmB4ltAIslbCQ3S9Q2e9
e5f4PN3vIAKCfRoOFwM80CaRaIuGSFzTatgRFDeef5O6JjRiA6ShIfTnD3da7lZGQ/+0asvbi9U1
HYPplP9ItHUkVGmN7lA7+C/yb/GW0aXIYLsU/FsqQOBEolSPBfKGCPUF6PxPY1k0pm4T8OtO6jnx
SrU+tS1886yGxkywkeCynju90DmQBAbFg1rt7CpZgoAf2WJcF+P9LJxehSLV8wKDoRosDksCqVMo
0pwedVN7paG8sCzld3Bc1ERGT0KrXBpdhwDrkFnjaCfEWPEHWPWzfHE7Z4h8VsDJG0U651jkw13C
usTg5+a/3NZ7JTH7IKo1feYkX3YbOtY8n7jtYnb642DOiqQrrbeGLyRZDmlEf37lb1N5H9c081aT
NaJqgElBbSt19+bVGM+oiiGWMTjvJN3rqhKaCPVgs9uwMialSkP8TvK0FDjju863qpYPwUeg7IWd
ofzixC8zx5mHkS93yYgsuHoqGYPj29qRFljjxgQvdMg6/pQjg6T4utjQt8b8y8bMnJWZptWVLjv3
YEJHY119hVKQ1r7ypp3Q+VW+7FLNVAxqwE0DZ2YDC4QMZoZoOcPs5nSonkjkZ/t8+yq+hI/JD0oQ
hGginD3E7i7GPbkqrTdwXI4gS6GmHJQ6mmFAPTlUjzZ4SuqugJIR71ZAHfBTJcYixm6p+RVWglCx
jVBDBe6Cy3wbJzlBBsH4cTrNlq0jq2PC3LHx8A78ATSyyZRYZrnlF0N86FjApAVMaXQbXNmhL1uF
qzMd0Mdcf9dW4tTYsE/KwLS6Yg+CgpaDiIMv9ZJ/fmVI6C/fofMSkDdrXO8+qYqlTN9zbDWUA2pr
5HZrC8v/Gvq7SyXVdBedjXm9zwk4thWEH8Op7HVYMl39cBZIpFUcb+XZmetc7wEBZTvX5Xe7jSCC
zLy5xRR3eKtS63LQ31HEhfS/LaKs1bE+9VBpWmGDdo5J77IW2cWBICsmJpF0lOE6iOJZN6tnxIlZ
t3yhpMVDYVOkdMvtsB8S2Yvzhshj37RicOnwkwqplCPm/qvh60pImxQ2xdE1rMEhtWADQYvA+q6L
ijXlPHY71ohOJXlePMuaUfS91u6NdduzfndqT9LfSqBc+lTlAY/Z/VW/ahF4/lrVf9zs438ODMAa
PDeZ3OwsgE2sptkQMZ678SlNHqkpg31lIl8mHaDoPk1gXL1ND+K15YadAKhlpmI2PzvCNA8jPPTW
bng8poMe5DA6WuVOstcZpxLOB5G8BL8PU7L/Hlasq8rRYvrf2FOTSzi4huxwK+9bc4FQmcFCqF49
Nhc9xX8WlBrSi/uSmpAKc9invLuULr9bBJHCACzCyTL3lsBKqlvc1Ls9Uk3Mir4EsWTl1bHkxgRK
dLbyhzq2Hy1wYjCCQ/dx/POdCQlDRIaYlwCP3JHWWj/q+KPJPGAjeouNOAtySszFOQMgzB7vrI8Z
wi8dbOm7zMn2ct4GRPY9l2cfMNUUs0FG4o1JWq7hhCgZ/pAVgt1oYj2W8WuXu+mfWQzujqCuc3Z6
X+M1b+FLy+Yec26Tho4KmG33ZhOXed+Idm8rx38TkJTwFIhksKqx74OzwcJOl4RCitpkjP54vr62
1y2njRhDDwoU5L/o142DLJRcN63kQuAnKmWWlQn9AkhvvLzWumKt30Ym2rsBfqoMrT4DcEy/+MLP
FoeZqr5txkJxadk09jRDOZHiMA8L211LqbicxGZvCQaHSUe2BnoVruWpGtpK3qS2TDm+uxv+0uSV
ZTPZ3Ta8izrTAIt/gBLt2YfPPpHhWmEpZWxnihZ3sdirSGCY4Uy/g/OE+KWkx3ErYeuLzt0zk6C7
/IKYid3Uq7XIXmNylHfqkqu2fqdEyVvgoBY0wKmgzvMwj4RTLPPwBRl1uCWojxNgL1GnQbPUwoww
JJ1f0/clLi2jLqOd0Pp/dYdMYS5n+Gc7oMTok7pPrMNkvrZRAXfTA0off0+ZjOatU/vJ6nVz10Ks
DDgf1Q57oYlLELTojkZscjyXyVqxrPqXow7R8r9KPUV9ULH2r6/Ttix6LOlPkp8c+gwKHjnm0b+Z
i4tSBoOKZSJ0Y68+anU2O80qH/y1vL8eocoO8O7fvfELl69Sf01bAAlfX8btP/+GLDz1izMq6u2U
PtF2DhVMZkrMCISwlnOFbGcxEohH9z5d1uQ0zuDYZwGReyxokhGxVMly+u6OePz0mbEhHMywF3ry
zXYwjfDkhyaybWqG1+URwJTgg9urdP2TjTlbXN5lQn/ZRHj5aOJCrz63jq+d8OeIBHiJVPbGdbXh
vJBDiPxBnAoNRqc3daWnj7B78K1CZKaQX5Ouu+1VLd8c48vB3DBlgHjyc9trE10ZdZ2/f3LsgRsa
2crKYGAFzQnIUJMSpLc9aSTBInuwl7kA/u22gf3JAiVFVn64e4BjgEPwXLyZNQZHTNizu3Z/WK0q
wdwKyZFHQXByLGtm0EFJ3/C/br8pBrpgsOQBZLhUb4hknS660qa6Ay8JV+u0OAE4LrqBC+yaEywc
wPuZthvIRUiszGrv6PLCebKcOmpHUbcNyC56/qJ+yN7JLluIjoH6CiEjIGrEXYAes13fI0zRo/lM
etMM7UIriMeoVobdmDQX5Pm2PcQtHINbzWkGRLn2qsEHl6pOPkTgMEDZ0K4sCdycNN6vau+u7tQn
S1UdrXu9rlfRzQNHNo1QF1/knbqKKqQchCm1vHkdgG/E55Pth/CpOJriea3sXKVIxnxC3WF07Jxj
LKJ+Z22nXXk/ub4VNi+LKmwUmY+fogxToGCkdsduEuftFuY9h8yC0FpS2hWNgC3yXIzkW2HpQ85+
X4nj1azQ/rLBFYoDg+9OwyH243rPHKQgMw/wqt6rXjt7RO3jrRy+gLKQZRNq3CUYQAv2AtCAkIo+
T1s8emqUfH/g9mY2DZUlQ0N8OmivPimL+hjeW58j8MUZJUG1gi5quJNJLxKjv6S07t3Z/XdxwwWK
xPEPOPFo7ArdJ8/wLxdcMz6hnzv/vwg4bL9+UlfF2T88TX2skwFF90Vo4DTNC6bdEYMVjMYXZCGX
AtlB1NOA09wl5GJDjEan/3iJQVGJnO2pHAOWc/rz21HhICS+afRxNqVyES3vynMJZfjJAtcjGvCe
cEobYDhMN+GhL8otH7x1MULjIUDpDVFefc6DjTjcfmfeGyvBJpOgpYljZWTYVVQQ6lL9lT/7Dc/G
4U2ApZZAQpZ06Uwu78/IQRN6+M7ra04Eeo+RL5WjQT3oQLzDonM+FeswJ/IDKn1HYn3eTp+gy4F6
PENTRuM/C00oKMmpay/0IR2mnCbAcSgVnuj9LeRJp4krgO2Xd2+3DHn3A2KAPn5zVjvXwr+gGrOw
AU4QJcEyeu1OglLqdUXwIqH3R0YbER6YKnYkM8D5c9M5lx30wcN3rBsWNy1hsavtqYtZtWoQW82h
t12o50OBXo8SljAG/5IOmmrgvLXbxHafhutWNv/etRJ5VX/f3EcWXBFUkEZELTAVG0edRAb8hIV1
CJFhQMtyh5uLFrxBNhNvZcgjIOoFFTc4XzIo3CZxs7hYW3Px+cmgg90S96L4Gm7Pf7Cr7qUBeKgh
ybxePS8Wn6SwJR/IAVp6Wo2kgxctGLhjSh0ui9RE53ZZyVY7M/y5ZmS2w2x0t8CjomOVxyWVvgZQ
RArIXhTpcmwbabxRKNAJwZlxIFN8B9XOzkmm5B01j/HxI/RaaIjY8Pclv8wefiXe5UzTnQtV63Vn
/Zn3dc6kjIOm1ZPesv2B8XcGBSN9/gjfVUXHiA9H9Oj+lZK0jrcjfsqGvILwJcCdOvAE1+v5/TDH
6grx5f2LOOVcuGmrXJ//d97Z2ztPVmDW2AqjvL23urrSk1O7BXl0VB9qjQRZ4Rqs6iwceb+B7QLj
kgYchJ08kc4/6BE0UL2Tak3XfxoJa/S5gKTf8OmB/SRH+7u7XBsK2yVnszVjd8xP9xwb1ZnZO8Du
OdmhLTdzmHTw7EaMEogppO+d8wMSz4NmqDHyoLuAgGcpHsVPWKH3KhWzfc+xAMAf1eBrTWly1Duf
R/PXuhtvb3SKkMTBChmV+Rj4PTnGxP5KomMvcuf2BAL+RuZmuaFra0Twn0g3/WqIJGjM8e4Wnl8r
Czi3u5n4VPPgznm/YJC2rnflDRUuo/u2xclPUl6CLa5I0eG18MMNGnUSH3qsurvx9/XraI5wO4LW
OQmUKyWsaS8xnyBMP4rvBNq/sKIk/xZIVNTPoaxgGJ3z4m4985xx7z1xK9f008mwstpgBDi/yAxJ
1HiyZjUWEhmFaBgfSsapsMdZBisE00d2w1A/vtMLwKCH/50Sf52tDMWKtue1L8yBwKIASG67Z3E5
KWY3TAcOpiIpMicksBBymaHrW5vpdPmjDN6JNyKeq9EsE4cL82Ko0qX0xe4XWA0SlIXq8Q8bHUQU
CzwSN9xzj+kAJdlRli5yoVDWhpg+/gUKkGKGFiHUHqddstXsw6wvgKqcLcYLN8BOzmhQmQQ2q93l
y/I3ZWJGLw/v7yj2GRgTSirdz87nQ/55fwHI2oLNFUkeTbGRQw0XjqiPNLvdbwNKgtaSIsDPAg7n
jrxq2L+cG9a0SatxTRQMQ0B0Ad/T46Ej1jxpGX4gFtwOP8+ysiLBa6IC28Dr2PbgJKzlkndr40Kt
p6NyJZ1D6lXb3/9+08C3FAR0ABJlgPvOghEXFiFqh/9OaTnK2ZAItVpKoCrSQD1x7mwVE9tKOqCm
o4QfPbNLnT36Fb3GpAAOhZnXXSgG6HEsH4pFdm6CiT5YC9bPQaaZq+IuEbr9KuXQ1dfdCRlRqXXk
G/dzgLudHID9DmoqpzZrAlS+3V5AXQiOmIG873jaCwZhBc7C/S9SCCKoV2oj+hJpDMMF3SbThO9S
0zEaWjv2SFcpOUlfFrbDpH1lA4zlZb5Fq9hTBe5zU7a+7JRRCZBy3IvVDQhBSOnAeN7IsBUTkWJu
Dn6KzOnMuW+kKhLEkZ1Q+USziK2VM35Da60U3hFLtHLvI+O2GheLfhh/ghNQgJjyIox1oeKLZYF7
j3UbnE0aGaiWTMFopDjJ5mASja6jGIYcFnwaSl63Z0PNey75PEJaoIWYHvxWWjr0c6ZLw4rZFM+U
OW8iCA3ESqMNlVfnv9FyIC5DfHmRjWxhAR1cJODuRlbLbNoQVohTylcm7wPMbPFz4nruBV0oAoyN
iaWHnX5614IRRu9u05XoVxzgOnTpydofzqzkqrkm/SY32HnBRRvDrEyTnZRTG3ZXZXxSNN0fmEBu
FA1LyRgRDOGS5JyRwZz00VjJ3eP60aWbUzz1m1a11xAWKHwBThC1pJS9I6at0bxL0kRlh2XrQAAq
fWBAwt1lzfGXFXLf2rRaTwnmXDGXfnq1IQZiWEIb2+RcxApbURadKQaIyHzRFp2Of5VOsHMvYiZe
X+/ZfYfqZouiXlOedL/dVPVoIBcFaasvzN4wh85+kCANI4uZpLWfsVPCcwJ6/CB7qGezLdD0V5X8
D38LYhj7Yl/uIZr3I0PoXMMsdx2rf++ZPccIhIP9HuGHQfSt9nq+xJxl0Sn4/MpR/Z0rWxOF9jEF
vUx9MXBg8tjRTb1YyoAXkRj/rUQglCghtzDKb92hc+Vy8kTaUk5+ykEl6+wOTX1p1/3U6ypHIcus
Z5YcV+kibRqOg0zYLl4maC7j1P9MhGEG5WRLgd4vOsS5+4gFxyukB4RBQ8EmkdOUnOGx8gc0RALv
v8BJ7849dH2vqyZZ8DqjBOIjasMghWV9eLYiQ6MBqCc07bCDyDH85nRQENi1XtBMb7QVbOTwJZa3
WVaKCOY/9nsbxVSaD7rddCAQ84b4ZhwZ4Wxvskf4y9IrbZ6JqnICZKC5f/8yOkbEahtTzmNgk/RX
H6jWZWw8xUQG1OptnVMpYDdiZGj6vAvpWWiNgRR7PmFMXJPu/ZLCF4cdSj8sWaPhvkcmxKOetkfk
bOWIl7WOaGclJEQrTxdOSdHsHpsQRN4uVNzs+dusbQNZt0HsPI4op0Rqug83WKSPMRwQcDUSaW+8
IRATLnGp9Tx0n2XBrB6ByrpnRzpeApAOOOMVwlQoeRtPasK7W5iNxik/Qu4pkQJnH+EMdqy86Kxh
H3qGvJD6aEToZP9hw4/C6x0EGPLzuypDptmGBsCFNCe3wy/vO6xYYNDKPHp6sYxsngn1pRbzjo6L
cIY4E+kRNt9iMSHT42U/sz+JR8tK/XxQ0h6RAo7R+5SDNphtxSyvo0vDTIyf2AgkGq1NV8LCQVxX
xxS+kWiUX+12QqB6KGJXLpmKdTUGn2ZtMFPjSp4tnvP7eTj1c5exZZ3h4LP+S6N5iujH4L35dnuk
RYBQMBL28axdRdHJ6ZP1ZxlxKW8yU82+/wNEe0PBwfq+4w1Spr4GGUxkuMB7/Iowcz0nNMaO2rX9
APaPSE2XpQauFF/zIwXTxHTlvyrDOQsDvKv1c6ecyS8RNcG20D/GbCSpcVM+UcsM/67S56yuZfZY
z5N+0pApC4Aa4xiJydwNjbZf1IxBkmsfLAUnnx7QJlAh5ydUNLCN4m2BM4b0YWzkY53tURFt09ar
5W8uGmo5DTuOvsDH+0sHUQPdPugA0pwewgY0Z3sbrnqCEt68nAW8Y3MVEtNOBHlWMn3Y1q4T/MS9
gWGydXIWLwWkhpSNOsWTzgLhxN/8mQA4D2d5zprmEelz3g97VigQO8sIWCZTDdAgGR1/jN+oJhxc
H2mhUzSNZpEpdkqTpOZre7Lgyl1snsK93PASck2ampa1P/GohlSVtr2RDcwMTVvwqb8+wATdx/n/
xk7wFCzdNjnzlk/Jni1f8PHTNz99nIpX7H78FLfAucl3mJg+SR5CC/3aMrXcPxYzr+fEXBVZYuPE
zojhmekU+0dKWeKMDOZ/lZj4yGahjHIofNZYHE2jYre71KMEeyiMRYVLU+4bgebQwcbz0QZDPTdC
C8CBErTbwiakJRWDCje0eGUFBVNbhbXTC3roTBOm9BLcudpLzFiJfoSjEruBSr2etfaZxd/ghX1H
HrbIr4/59Peh5Kwy0R9w/72btoHwT42Se43Ocz2yUZNw1i8+Uh56afstwdFtjFE7cPfVnRcRHbFx
v4f2Dmql7KGn2PNiPjjf8aLqjLo1g6u3pHVtyotPjKcO618Be69DZ28AAh9bhgZ7ICfTevbWgx3f
kym3pKaDfqpx6G1mZoEiYZ029H2ZJUCDee0bNCp5MWQowBvLLTmjYZtbzINV4oI73HLVnFixwGct
uqnBuvjEeBIaSrLsbMVZqrFrl39L1JT+Sqd89f3SoHTuAJJuAO++w1oeRApa9nQNpClELLngt/fV
FkSp/mW3pqMDlzjuqLbT3vy4h7XmTIh/9zLmx2D1MlwsdZCos3kc+MarRDSx3egDy1kwul0mV17n
Z93DY8ZYcfxUaTCU82SvbmuClX8y0vGJS0uKkWvy/2mV8RRwk/G1amMVGosyNOwdbj5EzzZDN2lU
BhnpsNAeGlsOO8ypNdD2hF40dAdat+shzXtBank3MbPule3trEkh3vqhRFEUhXhb2TzeOiqAkB9f
Nuq2Zg9iCbVZu9wuKXZmCh7MOeNfeboPIFlvjsXvIqEshkRICFrrhgFgEp9oXbP2vRn5u1mVmfXh
b+PCyMGRvIm492C4tS4HR43CMxp4BH8pnx/yUOxc2ArDFsPRXY3olfVCXoYLHH1Z+1nlulYqkkzE
OYoVfuLlQQ6pPcRryyfFNiOL/yySpNVX1+E4k2WDFIu4eexfMZxiILfMAcEgkaJzKY+gw5ZBI7rx
IBV1raq6ZMHDtLzLkwP45xunIwvkwL8JPkakAnsND5vfRdT0X7nAblZ/JOOgDcSRYOLFMtUDyHfH
T6V4aDQiSyy0MgzTcG+t4nYAcsI+Ud8M8SUu+Oxq6ZogtFgIM6DGpMMCmDERY7vp8hXbFn/2JIPz
bYcKopGwgIVw3MWdLqYNJjCKPDWt9cUX8UcJ/2TLSb52x6OCvhPirUqFtg+Zp7506y+QoBOOu+pp
qzCXFL2ndv9WnIHfLNdxx3JYUBuGU+1msFuqFpaWeUPF1/Ofk65MOJ0IWuv4lbwY9r58gTSa+kbj
xio6MLRJQTj2FAdOx/AEPX1r3k4Rri2n6vNShz0fR8ZOTavqLtOSdJCvgC6mFYP2+pAtUP8Yqgvz
Raqr0tPWJ3UCvABMit2MjPTRi3ckE1cLZTqfYU8fgqC1m/k6AkOaq5zwhD0bBJHsbeCUUpTHN6QM
YRSmr7J0wpgkTMAWAPxgQJZNIAL/5LXl/oZBB2eQdqID5zX+AQYRyeUrESaLK5pEtgzv+KvhR+3m
UfCfGMmVBcaccZ7qUUKFyEUVPEKSqu5lyHubAm5x3gPJRUuebH1t63R5nwfLtvcp62GBvIPmr2pC
jwgCp/L4R+V/B9v8zCjHVBcJv6/Ag/ZkIMQ5/obEKHzNBL5Z1RbirDedRSwSZtv1r7qxigEno3AQ
rKAhIva3XTk/NvuO2OpITr++Xw7yX3KJm05GZ28hdbdF/i3UATu/0MUUzQHnMXL61wjQ4ZywK+Q3
J4gt+hyZ8YO+gJSJBgiCsAw5mU6mCj6f2F8b5w2NE11Pos1AhIvplVz8CZfl5D+uIC08lrbgljXW
rcFrc1GkY9Y+OCSomueEJCHl3816jhJKpc/OR0Eok8LKTE3vSCt9qVK9Z8YENINJ28IM9EBGFcJU
gPDRWK6LKF5pXjqY3iq04DAilPB8f9f0MEryMFx6oxaOQDpj7KCxeO3bhB206H1F0nm1k9iWP51S
TvwHn9lO0ETijYpXBx+DEQnVTYQo/psv54KOEr9f6VUUpOKO51S8UJV5KgufFWnUWyj1XAnwKkWR
V4nttCXBMt71fbD1FiVNXz5YtcO/isO5gLM1TumuWFmiQAujUB2zJncj0lXLHdn0MaX8rzqGkslt
pjwLsXo4sArqw90YEnGHF5a+A3YnGMWsRGSd5L8UNWUAsoYLRJW3w3IQ/rOUJBa8ERWhYn3EIQc1
UcSKCl3QC27dqT3jLEeTgL4xxekWfS5QgN4Hb8i+X60XRKf3nYzKxi24KC/j2SK9ljjhXGTFqNU5
CvM/lstVnYHjhQOyg45lpCEtJgW799+sVUiYrh0wYBE76R4vx9XhPxFQVNkqVCR0wfW3wwJbceNH
+oPxIEBpdmLsTQDkwuCe/h6Umrhjc3qg8+DX/n1E8Yd++/Lnca92BhHT9N+G6SSIM8Ezj0+/+VxP
J2/df4xjqwhnFLhdIOzVgJ+2Lgm2iM9tt0vta/JdLubYG47rOyFLbl68TWtx875UvB759r/NP4T+
jC7CyTsFF0HV+lCX2boMVtOwjDb8C0YtYzyfTfkzBRtp9rJztTTiU18+qSHugWd/7q9OqDD3T4+V
9nOti62tuu5im6pCsUgm4EwgTw3DAmvC5isGgFVvv2LpczaODQiNL+3KdQT0cHWapidCi4mRuKDk
gx/M3Eyku6f0hwrHGdFvAVHQ3OBff11SJ2E1vJBVO7EDgn9Vx4uxhSF98Ju9Tu2GFPQ3c33YnrTw
FErvfpdAajWxlX1yNcpLRtzcd8JPa1SZkeowg5WZ4I9n2k6JlShF6cp0qEC49V1hGJli/U+Qj9cm
XAntCgkYBRx3BZ/Pz9+pyrdY+Ej8oxC0fzuI7kgWf87r5Hd3yHEZHAO9zyp7EUP8fOS5aEdctoCp
HRGsWRPIwG/CqpaZwSNc5YnGyUPFRzb5ANUE/UpjgtkRCB/QCjQZavr69J89i2QrzhXMQS/IlP3U
w8Hnllh+lH2tXM1VBs0AN+QL3VGLRpKW0SpmZUVkfZiMol8h5flUB94fAHG1H/ECWxHFLz0+ZPiS
73k9RvnnzfY5XBokEc8dU+RlF5UOvxiC0zLeaQg2UbjxdILJ0JAgn0x5+2S05I+Namkc2cLSyKEV
Z3QZO2HNB5+Ri1Dha9+DTVqo/yeiTPNe9ItAgfAYaGjfWBQn/4806s+gvmm7VZN5YheVZ/e9HrfD
safB/tKmrKFaQ3V2rzt3vss123iaK678okX0v5ituO83maCVmd7o6L3j6EfsDPgKI74i4bIPa7o8
9WbLq/j0pCCFe+sGxBDT8HxKIS3F4EAfS0KwMZLlnOi4tJOY3ATKaytjeg3Px3qh1yG0okNxvKAV
tVXgsvYDR2w8gvWwQEmJ+OwVABMV1hKRyN69WuObFJD938GEerSnyx84oau7F6IMBZn1HKVGTNW1
lPcuRPW35Meeqn0o/szpMA2I7tOMmJ0TiGtlWljLKhwxzTVvfvPht2ReHDJkD2ZJ47l5qszY5o4D
SwH7B4E3tMP7KnJwDWpsKmXNLkusrmLfVaPqGCsTq0MsVFLCIRM/RxHAHFRuXFALRct72/5jD2ti
INeKe1tzXFZ4gqLjEsUXFQ0Ag6dQaXnWBb2JNeWN/OLx8d0ssClO+sC0aDSSx8shfiD2YZy1G9PT
O2WHHnXgCg355VruAUfLeHvFyLC865RGFPK7oteyA7UDx3JSis7Pkx7rVZrHbNEwErympVemEzz4
oveJkvDlvvCMMw3d9qtPJIqkteF3o3NW8HM2aRmDZOgriSOMQ4yK9MXoC535efP4ZxPpdDdn3/QD
TVNVgjFA90H1AZ3bwpr8QsWfyUNPR/iGrqolUm5UA1wke8fCK3mARz8Bz1ssmbgJJ2WFcfjhfeey
L3XVd4ru9F6wZGCnZwPo4g/Art81RMJWwYNmSwCzlZtcxHWTI3VAebLMu3dUU3a0efXW+N3xMUhW
9IY9aMHSHsUFt0zQaPxzhwH0Pv0VNoNlJKQ4Kezpfj4KsEIrfXgCpK9whE5PDL7QPz2isuHArA2J
M2E8tz6trYz9o6vyQpr7Y1EzsZlULAfGjziUpHaXt44JJ4/0wjI8oHXXuDqoSBN90yQ7b1wu7WWq
wSBGwR7SpFAlnQi3/xj9Zedf36fTDdhkOL7QufpZFr/h7akdMrO83uyg3XhE2yjnncaulAUmoi0k
m8Pr5kMGzy2bCRn2ptI7wrmE6I6abCtw40W1v8jaCCD3BEijWKyt57X62biz7oUOb3K8D0RGSOXa
+3s4CMChwccL9Gw77zHvMeblfrFHzjGPgLwFoVEUEL3216nZCa8XIfbj1MzujlxpgBVleAsGbdvV
HXyAqWUjDzy6FhjePVASVQKTtrvGCtBvJzbMZBtPkaoZfNPVq6D0/NwuV1G6cXq0xBiRO8B6CfgW
hmWi6Q4vaKMUwqDLNTsXdIYM7iOkXY20oIwpgZPSBDbx70LoITIjAPViQN6+ifNr+/C83iPv+Je5
pXeRntEky7e4rMzbpPVdlCehuHz2pOyJmOk1gOR82paV9sLj5/mDJZfW07rX7/pY4qzJnmYvGVo0
A+79uR6qNZFi4YX0qgwP0YO0QxWVAtJSl8RB1Oe6vADWUASe6fO6gdjie9qV+GU2qOuzQrM+rwsQ
8ZwmjQnnEsW52HqVlNuKGRbSTRmQn3U16SCZifPCQgEZiqg3BmSq+6Qe/cppGiw0qBaTPQRPBDff
2sBgqRA4ehqHWxFIelQahy8yV5tplKO+bzriCH+rKQ+11VbwkGvVcyHaEk4yvRxEzBw8tXOqAG/I
WN3FVCfKuyOeOoC3ea7bOOrBj0eje+z/x4P9Q/YeVOGb/d2PrdEn+WkyIfmQrA8IPY0VOIrUOMqi
/yUjA/7yASk0JkWtHjkRIEx3VAkW+Jc4Xlak9acYgmjtsr/BDbLx4PoqErbBt+gQL0u9ZSM+a+Ff
NFCMJaRVI5OPRnzHkU13Y1Dvs8xClxgUO8vktQ7yLKmFlDFYooZBq7e84eaZYDjMkf042MMZtnAG
RTyyaNXcV4bmqdWYkslgC+iEZeaQOs1R7MMuDBUzy08CWM13K8isNzNUFevDCjLnbZ6plk0hdNiT
0Y7k+2ZXKNRe57FdKWeSICZFcEp5qrINxIypWWhCnyQPqYo/ZjDdm2SY1vxFcsUjKvL5+zwdlDCB
vrczN4g2Qj4vxggTL5tmpILoUAHwUK0xDbl2elyZsttiScShQNbU0VRXSYb5hwCBQ40qTyeniU/K
vNgd2KuYfys/pOQhIz4EaeIIchAsTWB2BEwufHmRuUNAH7/Sga+F8O7x+udm5ABsyx+FNDzptfBh
cgIhJ34jhhlGUd6LZoCwS5i7z6fNmb0tAhoXbXZ+0AhwnGvw5b4mYkfzSouaPvfldHcQOU4bUcrm
fl5sYsp1CaFtss4+SDbFceQWIHl7oYwlA1xdQmbJznAzuNBGBCXAiruDeuMLwunPg3EKa/v004lQ
ZLjfFxfO2Gqutynqm/HNCA+hRu0CqMRYSn1eGI8uaU7E7blCTe8JLbV4+t4JfQJBC3vTXFrc4NP/
5KorZIU5uu+Xx9199TBp9Oi14tTPP0Je7vl+JOf2gdw1/t3vbpPyOX9t4Spz4yIfhJt3DRXoMbzb
qIC03dItKWdGZDnGO1NhXnpS3IT4AQQ6Kra265AD/i0rxazZJU0B3lOFIG5qfCQUmYXLKWlR6YSM
srH3TGCkwXjcDhdP6EZeJCuFTYOgBFmtT0IxcBuOXMYVEjOLfBvZb8pmUhIHoasLAia95qNoPuG6
2YmxJ0G1ktBtcR8/blhYS5RH5I8wR4ALDRkpDjXl+JLVp0LN4K/xeHwyywdkqxDecpy+86pDaVxN
sebDJbT8lYxu6CadL7KNubR4KFoaDW3NcFWQGsn48jmml+xjT2Wq2AgDQvToHnvAB1MxcFj+Oz/P
qypuek+tcOUSLfcPkGUBq3qZ0g7ZzTZFHoPq7MRbV4VA4rBwxbcpV3GrCKx/thtFrX+0vMHX7MgH
RLiZw5FWlPnjXCEt5UaZyp6f26Zss/n4PZqQWggik/8699r0x4sWdyp/PgyCUL5aPe5XzBh3WKkG
x6gnEhUtrLdf19OS+tabWgoN2Nh6whmmMJlVZ2yoTqymxfvAWz1NkYLbqM+a3Bd8HumtALEpdAQL
PUT+Nmftw5rWzATIZE1Kc3b9T8xgFh2XQXCx5YyY/lTnWjCk6RcfrdIZc5/009qb1MSHODRlXs7N
GH1u6iHODHn0E9C1QsORNAND1w7dLdzn2oX5TJqqPWEN1WNGpWPsZb+Y+qM7lU7HxiolOtazLLuH
wVqkgqbseCmMgz3UYryR7V4SnkCRVizc1ZXKliM8JlhOxhA4S2tb7N6yw4b3D5ViM9EQX9g1Liwq
KYM2HQ0gPVw1V1eBmSevwOSz30DYHajqCM4VBzj+PgIadM8TrMgrfMtSwi8ovwlAaflwaLijQihm
vi1oklxiy7cRGpgOur0Z4wE2kW9aKIxQLdR3wYKOfw8RfKc+0yayFLOigqOnqsnk5Z3QinLuebLb
/uzTp87ld4HqoPupNBh+i8SkveX0N/6edGrTgBNPZcYa2z7HddWu1oT4daJ86yIFL8kD24x1nkHv
WzV3/bfSKwmOznJPvSb8dv//ZXVnjTADItwTxVLRqWh2dl2O0VsJvh33DGheu0TppFEQaK8nBi0s
J/tvkUkA49TC5psFo1uLctSQxLQamZ+8PFZezeVnu/2fir8ERyy/uFN2SRIh9WEBmXkX/jLAM/BR
PtE9EDBE7QgNYtONexxDLvCs0pthO/ehFmPT5hjSaw+Ai3hvfGnY1VURdl+zUEh2zeBsdclh7biP
sLxZK+VZDJQK/fyMd9utXEPFhEv2y2yJmcYvcHoNOR3TKC+i81Jj1VAlzqrBovCdD/64BPuEF9CE
Tzd5K7otTG1Zg9xfiWZuhFXDXtgKLW0ApVaVWtf7b1l82NE2s2LrrgujnUPdwx8naaSsEttR/tKO
V/dqOoFLc9RRSHFY0vfRlW5vSpskr7Kneqhmpt7FNqR6mEsEnrYjyrW05lnhaT5PpBCW3oZhUB8h
ZyDmo5Ygr98tkI43H832Ks3LW9WMT8IxO9/fDt0H21KI1mdXdgySwrAVwD1HT0ia28NbVcdeZDu4
aOKhXgHqrnbF+0RqiwYMbPx583y5az9ikgPD5JK7LnNvMwRlpjSMBznIH5P3BmNNM0nGrFVvHI/e
DX8KmnYNq/UFUnNx+VHeDPg5GaulqUwqencMBDvFfrCZW8+ETw6d1pGkq1fkuVXWPZItEZ0R817H
6Zv/8+BdoUX0SnY9UU8z7WeSX74j7SHh3Mk3T0/L4N0WXSINOh1d7Db3JQ+6U9DDXkwynu3OZPrV
6Mq4CL+v8y0j3TXLGq8S3C0daouQLO5QiU3PxdBnolZXyCKD2N4bkCCgiCrAg9TDFbHs/FPM0wse
HrzS8xs/wwwOkoTRmsBB8dOkmso6djKG3nfS0hVdnY4A2jCWV8k3UBFgxf+b9w+MLwdn5yF/2ANG
N4cl+MOvSB2GxoLYCFN78mhPmZRX0FMudWXgJnzUtWccDMXIG6QoAS8O7X8gpXHmy/tG94FUlesO
bHF5A1BLyobhQ1KmBugTH+utHuvCGqJOk3WxC2Ern97if52Hm17vJZ1a2h3fqWPwUnpcBOwlK6VJ
OzkmNzNeUQQBWKIvIbwj+ZV7VlWs7nhMTQaOeN7fR+eiEwG/5K7WeMlZSogXj7PEplM/2MNWHd8Q
V0nCJmQW1+xqkEYct3S4LDzwDSYUayYG1YmMLNY+0lChmYVLGr3huznZnGB2peic19iBLE3m3ogJ
nTzklIeBUjKSIR1ou/g/SOd8zqlnDd4rev7bywk2DJgieLRHqMBOLMgPoQtFJldAyEWdui7Ut2SE
yoEyIjiStIZTyf7VjY8iQFytRZjKps8/6IQpIdLHI2Rq8xJTA1C/dMkkQGGdqPql5bfUaf6kcoJm
vwSCR1mlgAvjJOWtb+Lo4+u9MuTemt+uxrUDD4GX1qhF5Ji/SbHeLengdMJ03d7oM2bbC4K8ir/V
gVfsxUmkB4n3BiZONd5wuvX54BEHwck+scRBqEMnISjRw7tt61d1yagl7mxrziC3lVDYeuw8BDhs
s3vNxte/yPmfvpPrGURlMlM8alKsHC3mDT0xmTWph8BTWDW1lWMXhvAlph7raSnHQoKIJKQHbPkc
f7PHY1b4ahER4IfSgv1PffWp2RZWWTS7nnYtRdB1vgQy+1e/AZgoAH9yrs1puD4Z+NXfvIFjagN+
rbs7G1xkZ6WLtDNVi+aBsWfo4DpfDKirGIhuJqhZSc5WgFYy5dBy19DMUdcLxmVT6GuBUFMBRIx+
KzHgAgTDbrZHiMaFCkm2JqX5LCqh7l4lv9Fx45p16O3DfTraIfsCogXgj0JUslqRxy0fAWFyKA62
Nm3OeT8xcsO6YAffyDDIiBRD9I4sClJ5fSleqMHZnYdDhSenOtOwqwrtJjFHXjvCjrByAWXz97tU
JmmZan6oaiTdFaYCNWWQE7gPzyahYMH02iKi+aTDek9b/wyTotXwQVc14Mpf3VdS+Xz0CmrmyEGT
B5P3LD4/FnUXdyO/4ZvtkKnRTDQhKf2kBHhp8mvdhYq0ctg+S/VuWp5bzgYM+fC+9C8T++hRWciw
OOE6vzI5KzS66Yy3ngx0e2qm0w7qin7MHBbCdWgaCvMiwgn/fJ2gf7jmCkggUJzfuojA/TQB+4dF
NeJPYC3mroc7HlC0xhlhf599YD4PoZuH2oO3Yf+J8WAC8EhIp0QPsDX2z8oy7qEedf3Bq/NlZxF/
GR6TL9iYGLC2hqYVn9YliFSU5NQSBXNg/0l//l2g724qrucbdt4qgP0Cw+x+OQdxirI9U50vw/eR
Kn9EvWoAdHWzIVyK8Sx/J8kGEq16QsLTfrI6kjmsugcCtDzeMzuMDD5WQAINbu53LfsLlAURe4J/
StxINWP+pE7n8ugkyyoQQo2m4T1gs+8ttpasaSYTI7wfoSfs9esIS+/Dt1P655dUBcH5dyLn91gV
iWdGbdytbrfeY63FT5eqaeDS9QZqEqk6zEi8OStj5ydNklC7Qye1cRvsu2dHCcUn0L83ctTXU8QY
fhqlvZ5cSWehbh5RlhLWei5GW0yk37HiJYJzcPgwxxv50IWYny53dTmO3EcJVQoy2LETU2pwCnZO
oOAySazBETQavpB+BMFrwe/lqXBGr8LnfC1ZEUJ8OcnKBU4hmsmUur+8she76260pFVhqgLPD/H5
RV9oj9WYgpjRh3p3ycUhyH/oIlmwszDYshKVWXrcJQ6ktvrB9lKusqsDOLEUYASGFY9sNTbscQOz
5hIQ6R0oPIOoUSQU/lWD8bC4chtL6pVnq4B280krmnwRcvQWNxPSHnBLR0gq6fyNFsq4ys3Vvy87
xlyDSMLQUaoHeeh8YmUzAMnJg/tzlNHHvEn9hCRWaobXh/Kaq60SW/fpmYfeV0KHMFIwWPughTvH
8cPjVEevitiCN4NV7YSAWdvsk2wU393NUPk4c9D3ll9rqOGvNU1QiC9/InDBhdCSPS/MZTzfPGih
KVMp43/7MxEnujtIWWm7FZzzc0BJfpp8MjMDKgJXeYkA+1A9Ep2G9WqXD5us3RC7EOiiCJwMUKJZ
hbMPPZl+aprnt5jGwf8RRe7Pd/gobnCzit+PFw0R4uD9nywh9xa1ts6GjDBojdy5fQ/EGzwKjhcc
b9flARlJxLvyEueE7p+bJ0lx9ed8prS/6DUMrI8eIYNXfuhIv3rBYu+AGbll6TWwe+00CKYqw358
teZHl2H9jQTwjPDI3yqx1FSvoRYexKWB28ZKO1X4L+n6mBcNTsriBkgx7GRBRnuH40DLRgBRTjYs
ZS5wyvifFcJjOSyek16eHBI7m2egv5SuBgzQqt9ebJfJ5dz8vWz5HKJH2uBKejWd48/G43XgleZO
hgSvLj0RFk1a00pHw0jWYTTbeCVRlH2QmrOfAqy99td/3NvwG5hkoX5L21MIaYrN6aWwSn/2YWkA
sbPZ7GOiKB4/1o2kGQ4mV9pBRlY+ePf8u86AQPihq7WMxyfgpjedmkPH8ZwpDplVY0hairGe8qun
hQ7ZdR1MkJyoxvk+DSXFReQVrdAs5tDs2qPqs6DFRdZDIT+fyxeRu+biL1Y9zFcZBpcMxZ4cEFyH
F1X/HRH1d83l3TpV9ipXB2pqkEs7Xtd611hfLmAc61W1ZbUigs59/blOicH1pAdCYj7TuxzrHCsZ
/04yBYLYdfgr46YDFO/H6FDPLaJKCN8+aFI8gM1/fJlo1wKYtbBSG/se7Gg+ZYW7Rz9+yNUaga/+
V6rDXUAjXnfyEP1S+WLZgtA/sylVtfigPokH7Uha3ZOUHM3jFX0HkKVymgdOoHTjWrc7V6F/7ayl
kRsUsu0FJmuuiWGzEuQHOMlNj48E92fBVE0JqCHh3trmYrmVzvYVMTeMoq7dR7bTVrK6zMVIAwzA
niolHusoPJ8vdxdW69EhluR4O/WAWkmPj56Oj/eU2fmG8Z9FVkG/9zI1gXKJzyjviyBuN+cU5Si9
tdks05ni2OJohERlKIUTcnsJNWMBLU9MeJcSUfCpAVTqLI4amr8je+jSno6+B6EpZnwQJ46RdbNH
iAeJyMqIGMgD8+ZGQykA3k3/dNs2oR+GsSR2spSalQ/mr/PQ7D/Fpv0P433ay6aHq+vpqBopMytR
PzrKlO9F9aJGE91OTaLq9p7fbg6YMxn8r4/7N4SaR21t7Z546VFun300yjPRErdL5haOpsnWB+/G
fQtfMeMON/zSTJnEokapMEFsUT2tHBhvBsSVxgQk37rDkgWAlcOw5DrocIQqdS6JzrYWtRRkS3m6
eOZy559FiVIVrer4KrX5CGszTaJ7WfE0N6eV9sD8js3nB/Di2WK8gA4lMjC+I+zHMA5aeN9yh+Ku
0vLURh2WjeABrTntl5CSuszmSal+VOacw6iRbdN82HNkQYqo++qG2lFkeIidn7H1JFfv4gIjRBSQ
AiUdqzKNdv4HLqks1BwSTCTxloxVJg2FLliH0CbMJMZ+niPqOgAvMsCQk5CnChi8HZYQFj5mfHvM
1szUqGHcO7OFg6uWUdTXqsUM0IL/rzt7rHdCMhPzVHb3tAGLKvXxhGKJpvO7e/5bb8Kx0iZYeV7n
zTysiz6LVOXv44cmC0WwdDbvUI8dgj3uEKswNe03PJYnYuby/MAmz/0mAaxZYlNRFQ0Fb1rcabSg
ApAL808gYP60/CVbKYYj/7F3asHsmE5dSrD7Tt/RVLGEPNuTT3Y5UmbK/GxsakfVZL5JtetbaMIB
lH8J2ypohv+Lrb56tXy0nkhO6+sea9jEaoCkxiJ6GHROw/y17ap077YacrVD3VCQLP1NskyzO0We
dDrMgJ2uPRV4QTvLPrtOvcOeITwb+913tX6NcFwdT7w2Rc8D0NoX6WB4OWn3HkFgt9xT4pjryPrk
iht3EdIv3ZZS463tawi0R4TTMPkCJMJBgvRLr6XJbiX0DdBQl/qSHFj/yxqI4lClGAnnSh0IWtno
iSlJXekLq4JUkrC+nkL2VJVFJpdkgxaAyTte4NM1ln0slO1RHnObd9WgIRnwQIZrl6UlD7KAjKe7
+8FJc42fKl31vOIFe1C/SuMbME6R6RyyxAe+8ZVJydYmOnZUSwri0tWeeP94X1iLxSE9NryrPcia
vCP80FCfrHMcgasIMA1QJcQOuXS+XNvp3rjIm4yYFL5lqsgSsPPCmEyVLfm63CGRGw6ga54KM9dn
nK0GNdu+CnfsOOxmvUwEl5pcp2U25vRS1fEJP5t5zNLLWWoqkoIJKuGHvDAhB4E+JJpJYJu/7zEQ
/+iLtnk3H9DneFoI+qxX83JWWc3++o1S+V4RAj56NgyAbxvfZtZv0iNwGQMfWYoI2UTktEkhEIkS
b2NA08L5ZRZzk4RCDpxpllztCe3emNLYMy15tZ/KwcWnHI5wPV+aWJ28dUDeQFyRi/xc0RgW/YAE
whHofjj9mBns1JTMT9Y4tKbav1FXLZs5NaA668V1PDNfa9lssdD/7wTYMVnyNmFdWwhaygzPwod9
7tZiLohprYviorFFuQE4A++nC8sh0JkHGN2z2oD0NkKAtPca2g2Y+h9gXncSlCMoR5Rsmp6YO3DE
wo3Gcc3J6bDasABnjvYiDzRqi5kdA491cs8C4K6gokkIyt5DHoya/CvLO9IBo+yxw/GP1hNyViYM
1AGc+iyWrWTZ8maBE6whAriY/1Ds3bwVqkMHGDx2I4v6fA7v3E2ONf+A5fOJ8gTI2DW0NPhKiC1y
CwZp4YbjIcqlq53h610kfWxtjsRDASnijVmiAXKetRMtgXQ5bzMyvRDcTQ61HVNasx2P65D8+jtM
pxeNb3IXaMCbT6oydFa2pxwJQBEAy8Yn4BSqVhoxcWt3i8XaXR+XyWysvaNPdyA9sF2sRH5veEq5
vMJ19t+2uw9bG+gc2yMGN5jzNkHIOaqqpiQWWch9MZX6AUAXCIiUZL4MDts2G02laDDDAXBo4ye2
preeD0StO8Lxtr2EL5vHWMZSV60FK2+ZaiAcURtjLYgvIl08W1RuckpmzGsulwG/DNJtz832fGUe
KWTyIGEWq6ZWGERfOHvZfHGpRBzxj82HL0gH19JTh4RSSFKR5BCaUoUnjx+DClo2yAHWGUzauyqI
jHrh+vCs/xmxBx/76zSzXCyPD25sZyHyix+QLj2qPMGEkgbtDc0Xd6qicbJ7A9csV2rL/ESsxLNb
5jdU2G4bd0tDiCdFiMt/sCWVormjWZ2+rgyZSm7Qnbi0S9JlasFjWkU5wD0swDIISbLGgohvI5k+
MK0lBG+lFv0Z/Xhj+PbGOz8MxtAVMI0pwDVEwcWEGI4qlPj+d0cycQflJAACuTiQHR1R9oI6nRgi
/FUUNtjwAdlYKkvcH2oIBVwaG4zW9OYePXgyEVXwtWQkSgVUDFOEZKvfib8UW56/t1HJiJMxtXAz
4kt6ffRLDyXrZgT5ijma0/1AGWSgL+2oilGpWuI6quX3vq2vpF2KcabiU3UyWH122wrEZla9F6G4
MVSqJH1vhDlFNHQ513VkIlQmMsOic2uCrTGZqLGjobOrT1ABwLtwNLbv92kpxSecqxXSC01d2Hq0
/bsTSKjtxs2o4fYMmRsx2zX7aLAoADvS1oVHCRjYAauL6YuJauK5UcDo3MC9Irkd878qqb77gTYa
vC2P/SvhMTe5QQcSsEDUCgHO7fIZuS5ZkpGI/BJHD1sRNa10FAf4TpdFwqKlyxgPT9fANvTki+6s
mEY9QqqMRerzCCxjdjftQvo0OBZscXoiUqCybhdGpyZfT3vI3R/xoMxXfKFZgHdA+OGpQVlkf0TK
kM12EKnwBmub7JtWNkYa4sMnjRWfs06aW3veyTCzI6zlA05Ay0/R6nuH8jwEIfxu+JP1VW0KQ1XA
lfC+qV1XUK5ChLq7Dhcd/VDu2Yd5vzA5iYuk4Y5508VREehWNTcoS9t047di2LiYAwD0rpHc8PDS
1mn3PL5Bwsc2YlsI4wFg1qXq33Owp1KbSnL42mZa8i1gmRUPp+wzoxJ79cxgz3jvqluY1r9iEQB9
zR2UKK7qUiAhak94iQNaHsXdwUAnCLgkBykuMhTPmhRO0jGX8sVcMd+UzD+VnivdhTVjW6iB2Y6O
QCFenpUNsKJvHjFJTLA9ur4frD1JFHcGJfKzuaKdAuc0/hS1BLnoCYaQYpSxmMsCwyj2FdMwFt5p
2+A1XHSNo3yY6mE7zECFDruCMFDMVm5PCpqWgfrX6SI6DCLN9WYabUX0tBoduMlkPSKoa4oSgry/
kasLko3JChSP1Tcoe/oAsox6c7RPN9MBcSYZr27t9Vo5IUqYwNt+bYP5JX7zpeNrJNCntdrb9Ezk
DqrROSe2R0z+/pFusFDdbJBKHcBYb5w7GfSGWjAoHCBjhtPP7ojrPIVWmuEe9EerL9W3SZO3q3ie
1opaYUBXocuiLeLrclrgIPvopoCGECcDl1ABiyKJhyK4Y2PEfDbt1dolHDKl5O3nWAP4rrU8C3pK
+C8SM3xGLMbt73krFYgVWugC8NRS2z5As5gd8IpZG/P7L/neHZbhbhMq0IJoL1X8kICl0MXRrg6T
XUHd73KDddbTNyUM9k9crwxgvgLL5LmgtbIuvs+pf3xCInXV8nxsUE4o3vIpmLackPbMH0eoyMTs
M96hz1IA/70gcBX4jhchqO07BHHKO1GvTf21GXi1SLaiWEq+xvZB3EPVn2ohS5sYjMpKWx95s9g4
9qPZPsi/vazW0ytU6BScqb3hbDYO8IdOWnTA2AXhnUXtd+Lox+Tdv4O4Uy+Tx7hHBCZWzTQ2gxSx
9RFLn+VJ+t7uR859xAs1qDG61Y0yyZlT/LlOxiT7+/MKMFPOftz68BARs6M530nDPwIc1KInzrN9
FO2Qm6rGOVUyF9bctI7Aan07TyGJDOa1IC6XMVUBmpKq11BF1UMY3rFFsZsW47+y1Bf0FasclqBM
I+Jf7Ndf4I08h+X2ZsmeqvY5Beha7JyUA1/Ct93hKEWVW4X73oZkMyrWOP4Qj10l0mDLBwqWYnFN
ifz351VW1nEa74bCyOR+HO97X2mG5hqB1djJpvZYQKf+GMDmb/kyf8Gar1vbUPmMiTu3ICuBU4ec
MgyFMflKIzZ1T3IbR6fSXaY0GN0tobTwsH2zR6j3qrs+5YcVtx437QxP7oxWjfaGdaqIccQ09W2M
K2jDV46tszROf9Bu8rQjlkCGIZh3Y4uCAulGLjU2Hb1VHagDwvAhpmQ5PPIN9A8FJaxG5yV4Bigh
j+GmJyfw9ku7Jb8QBN+XA92upN/83pwGMoumzucJUAA6tuOVH3LBQ0wurZEG6NUZQNSUjqZ9lqyC
RlhMGJ+5Oi/+QINfhttwhL3QNWFUeoccHh7GdDdlktNhrYI29USO2qbDaOshYN92nM8ls5OL8EsM
CB4+jLq5573RarXEbcCEG85xn/DhxysA0lR9+Iab4iCtaepjpjYZp98c0FYMKdewwSfmPIVAYH0v
FmfWtagEQ46ZUKqMUMNZw7RHMu5M+4x2chjcBT6uGx9WgDrBQqFifVRCB8VsAAJ6gaZO9cmthnuE
+1KZPD8MtevFvUFiMtkooLtIyO0EY7ryslk5zAj0ShP5Qqv7Nslwzu6HI83A8aInuRwGFpqqsyLy
iEArt1hcPJaDKceTmYoldvvN4Wzhw+lza0Lf/OiOrAPrsGoUf7CxvqyiBV8QeqvtCbPs8FJxSaOz
vzrfenpF7swk4CCTTplUhCiz8Aj/BqfC8YmMey3GVVUrAAWmgTXomAdZlqZUwuU7PAinyGxWuKOK
1jQ5Z2KtpZvW7rhweo/p4a8G5XG//yeBVlwsM428hDfRFOnBB1nmZXSuhgwnwTwwAFmXhJg0b8s4
489ovyz274PYome/7c2DfBY8CQdgM7S0WryOAPztFrLvA9R2+h3pktUo6AJiONj4+tOyF3sJ+JOZ
Jb7upC7Znh8LtMc0Gjb1jRK3HGfjP4t/dDdzTMjB3KaYjdLLoGF6T6xGUw2W1MsmpiCDVM80wi5X
pjoEAWaIpieV0SgUho3+zlrtdmTDbLMj3U24Y0dDKqDrhlwq1ep4H2vo//w+jU8lXZmAw8ZbAfPB
9NVmf8umplvUCfnVaIftx/Xh/yyiA6+muDBu+MnX3WfGcfZ3uix1JnByQHM5h33cn1G8f/caZOjy
pi1ZsH6aJFg9elSsdxDtztRVuiNGyqX0UasFVi/DublK3NwoI+Qkk9pVYnN2kYvUct5Ud7UW2hTq
DWuckGTZy5jQKttykN9TQNNu83nBkY+Od1PLWlvjl17EQDLnnYUztkieILIvFwYf50iPvGQH28ZZ
U8YsE35Bpm7Cd29n5toqNVYG9FeKbQBd+8EbbC9yatHbwrIEB2I9k3zeQHQ1Tm9ZC2ZaViwk+Myp
q/AReuDRoF6qTmsnJ2Q9NZg8bdtmZ+Z2qzPD8XpEcBbFbNRfBD7JX44abB4IBZvnxaatM6/qmgll
YzPayBkUt1Fp39iwFV7l+GirTiHmRuWY2xmyYu9U9MG35QnSEL9QWY22tPoceXTze0RjzjT8vC99
NpZ4IBLItMGaFK48CQTE9mXQaSx5mVjg3iBqpGwR9RhO7ME0pyrEHQA2c991/bI+5GkfXrF7bbrm
l+pFBHe6gqNdDEpaZeLFUq4mqoO5nOEEc4oRoIl0NwgDKMgtjWWxDdQqaGDtJr43IscJOdU/NN9F
TK3l3eY5iSkVnEqcTJw/0gqmXLZHh7bRL8wUtaUid3zd2+L/eUowGyy32ZKz49E0N9mM5NLu7MYh
VpsJddLMKIcs04HN7t8kaxt8sDAkT42HHg+Uf8k92k+MUC6So8Rf5bOEjEZUZSHdmphJCJ7UbkoJ
0Co2MMhtbK8UHWIwZh3aesIVK71xikeM0VvwmzmrFZ8Lr5NeBTsCe3QwThgHa3rr86aHIZtjRZKO
2vQ029Jtj4jJXQV4BrqYvVHbC1y93nes3d+PMKVOjCiQ+8B9NQICLubCJSRq6QAVMFpupRFEwt/x
5aEr0LrFDnjJe+JJ7lr2J95hesQw9tmr8d/AKRudGGJEgTmNsOhJ2nX37u3HGKNfKgH6iRofg+7m
PAru6tldux2XBbPsJUsToxaGJKENAHUGjXdzmgKU5bgDQuv0H9yo4H6xCi1pspaCtMHaNJuxI4oA
vj7EWNgAnPFba8zD04oJE0sUnp4YCCDOwUU/DIBvy0/aikL4ZjsL/TJq+ym2UxpPhZMFl7jtsyYm
N5oZPL3OecMYFIpbhkbGb04NWzwVpYTqs8QkUjVShdtJ+UhA8gaZIm9RAxLiFbQeAeCvsuHn6IzQ
5StAIPIAIGFq8G9fF86JiXAtKzDV0TlmWOj0dbx1otXVPqF7v0JuSfeBH5aZo3Ruo9JClmN/mU7h
uDCKjsaQ6sD/B0aaMfh7a5LDhjbLpTe//T5BbBSPaJQTDu6tH0nIRWNd4c3CRb8s/fyohXHUBc74
l+1BSOLEmDHBDojWnEUgFwc4su1pZfRsoz91zbxOl1EjGhNA6b96of8RpZsQOJgr2l0B2QRj8nii
+yAJz+7DMktkmiHhlL0HmZXN7xDVJg7AzDDE4Btlz8rr+IfORAz1yrSbwD9CpPTZ1XeLxVPX6SVL
loNzKnI/CEwqtA7WqABQ+SL4g2owtGgeCAcBhF7mnLUKeOQyQERQ4iWst2S9JsMOPjRyFhNcnIY4
2NkWYR6cGF7SJMAexb4f+Ihv+upqYbw80ikfSwJV67G85cCBmm/9NZJ+bSPAuKqO6UJ52UorBLw+
ThFSg+wJfbkwlWbgW0+WXi+T0wI/NyZ0DOOCTAiQt0Ao4sbfCnvMOu0mH62BAGjJYCCNCy930jkk
mmnkwssx9PvlThOUe/tt9kxDykmtMrIkKck0iyB4BvYf9uyFRq32kGrHrJKtP3AwF0pR5bBoA4Gb
DY2BIPmfIlA1GUEV0HmLtiG+KFTls130OzT1vT3qhv/XtQREp9QN+mTgDhqZ/HIW5t2PfSPhm8Fw
wKWH+wfK45/CIPkaXkYtEgw9+JFUhQhuX/yf+6EH/cXD5bXDacsIN6s/5tH2WsePgLg/b3Tk56IP
w21tCKUU1q5Ki2FfqBYzcDEXV4PBVL/Q1uOsOL7nJq15fS1qukLuQGcyCZjM4+e5fzaZsyxOUgLG
PbK/NeZfSHYE3XQyqkFNLy/m6UnaDBOAoXIkZE7eher3TQBsmCqbVYVH4csQoHustF6xwnif6X92
nfsOtExuQhxNJR19zNbUHCYmnmdVnml/8PFFy0moLnFQs74hW9vDUly4Ct8Wl4UVUOdw+dNiVbPW
KhR8zz5t1LvsH1KjoyPNyTqoFPFp+JS/nVHeQFZvNzH8XHFfdp59S9Y+vgqY1A2i7pKG83nvz/Gg
zTL0PWXS+fsMRqsZETrTqN7IAvQOKxiS3Wl8D6tA5cmhwCnZcFgQ0iViFCgFMWHA+FiETlKVQ6fM
bLPVcFD1FLz+aF++0tbiS2Xc8QM1+waFFSwE6Wv1vSxHvtK8BH9CcYtoMQeOQpLlb4EinnlT1NTf
s8DWfLaMhdL/PyfZvXffwI6y9k7/TEP3Gzfw0q+i6fO8wV1VFA/L2YCHBmQ0PKm11RbUfAoLWJvh
n4vDNwP4zydwq5ViE0W81IhhFx5sD33vedn00e8PGIbNGl6STSlO0WF30IiOffVPLVvPywRP4Ia0
xegOi5BlfejvXoIUOentvX859gpiPZpoBUgrSHjoK7BGw+fdwbBl40YUToK7gxDHU97qXprr8nqE
EZXhmvA8IcerHwLqSjlpoLChTbwArNkQ28fdMgNJpyvtHxUVc3foNGj2Kx/iA4N9XIt8NF40BZz+
6/coEaM5A2Oag0NwpvFGDCg8qQB19S+dsc/nZETEXea4B4RnIEwruZ8ZF9bediocrw0dP5XREd1k
ovvTbrvUilTPJ6rIh/gEDi/QjZi7L+fyWuThlfs/aqNwLhHiSQtQw4MhGa4Aiw/58w/PnIIPazcm
G11bBiiRQHGLhdDkKcJIW+/9amLbAXY227EDhTvcJquxATjm5SjP9fIPRvwN/Q5KlRA3PcmEM1Hu
ocUOc1fM/xo/pq/fX38kjWMyMUXZb1BlEUAS6byCOjSxVEsqyJdoc2PsGBIbhviOZqkggWsiTNmd
YqPW6uuar7OSwSMxJPf3YVNnGNK5y2897MFIOE2yTvCXnJV5NtyM2kyV8dYdY3BVNiIHX6/vJ9Md
qd5U6zxqL8tW2dXLLUxaU/EW28Oi/548pdi4pu+Dw/YQCpLCLuPxuxmKBDHSdckuf12M5EKkq3/A
r5WziNtTjX+76j7J8bfURQ8+TNuWYwfjk3eJ3qC2Um2T6GSEbfKEnelGIyzFZctUU0opdrbN9v+F
BLycEx848CXpZeuAiEQqK/sXvxLry2CPXdBeZZoKmjWpom9E/9Tu90L97gJRNRZcg6/0f0yRsdob
sQFzzjR8vk7dZ8TkkIum6p7CMfx/j+KLxOQeGjpGuQLZRUjLSBiFFTnvBzbd79dBffN1kcfYsshE
wJuV8+c5JevJgxByaME8LRGBpDY6ik4PJLwjD8Ahuc9hjlQKxHox55zpRRVReTV6EBQjySVixTQo
mcU41vwU01Anv+BE80WFm2JYlSEkYUM3LkoU3Ku+Ut59ava97gUp1xJZqK/UEvOOr6gkEgF8ykee
hIbu3pqnzbtEvSAmQUz8W8cfDTegbEwqa5i5lbnPmwzBQizJ38JuED2CCIa7Kpt/ccvpgnPvD40d
270sxl2vj1M5l7DLUhCaBk6fTN+0vw2gdeaz92eTQFdlP24MJqVin/DmiLC2zwi7B9T2nON6Lylm
Vz1lkhHDiUaM9fb67D9enHijCOh3orfOgCEPYTQGVLXnsSoMYTMduMZ4vD5xKIaOnHaRQUUeLpbM
iX3XM71s5fK8vXC35bJ2YGxNNYXEqcm1BGyB/tZTdGeoAjeP0JX2NbN654U6ubFAb1aTjQUcjuhK
3WU8Dm8wfl3/k7Bg2ibG/hptfO2pr9k/Nb7gH8VF0wMeIzb+rtg3zfkye9b6q/EcSlNWMX8xI/ts
jOSivGRl+kNTtVCEk/cwDP3RlQfxT9tErSirfQNXpJLPIib0s/FUuNFP0AEaNCJw737WIAYFeiCR
AuUDQLxdl0mHBIENpWf8JkGV6hEoz4KMMVtDDmbA03KsaBOIENU8YTk1IQ9bn0Bo7J+ZooRE8qGe
R2/TcKNBdTnrNro9AVdrxYtKRh1x26HbhNlqWUknuZgGs72PNwJg0z3jYKOqTULmqGNITKGPAmLN
ByfiLhxZahHdayFa+IM+tiTMoelZ3OPqzjin2Ddvlk6riI+16ZQsAMVvq61mwMp/g15c3RFeBTHf
+PZv+zaNWkVNdQgCRbrwz4ivC4WPyPx2z5bBhkGrPofacHHJjgludsoFbeNx0h5wxEJ+1iaJLX7x
H87G+QTd9gnl0L7yYr0mWSHKkeCS+FIyAKdy36gkqOnvRf5OZZH/H5n+t7QrHiETcWI2Uw6gI2Bh
CGdlqN+8msBvST9pGa82hCulX6jfoVhqPj+K7/3xJN6Q4u+kju4gCxmsKypdR6FGLsHalA0GFpt/
Gs6pSjiW5saxyDyclgdz9gR4+YVBH0K/qDDlTIQqVRcuPqx/gGa0S4SrRYc4FUm14mxPDSevHbQt
kNp7uvn46nK1CgkMOJ6EeFz23eWusLyFvsODxfTPakMvEhoYHPW9Ufp92OupQhgm4U5aQxEJf2aW
LrZVMhxJMS1wQeBKLZQ86ZUAle+RBSGcdQolhJbJwUWFE+7+Xonkfp06Phv+JSqWhWhVa6s2IIWl
veQSo6iXGXMd70Ws8z8RrNd+GACuuxpqgYl0nS0XpUSMq1fPHkkA7omEeOIEnd66WzbqdSHRK4Nf
79PIG0BrIVG1XqTYFBcPLD2ACoAGppVxJVmL44u64Lq+CuzDNpH2t3XrpeB2RqB/JH59taKb1MxY
QhxdiKieYLmi+iCMQWYOf+RxGdywa4JoO2wpaByldbAUQsQ+2odLr5xq3ImDbt4WWuzQwuFIq48R
XtHjsfeEt8v09eTCupaTWpr4pLa/36lX4NVCDfLpbdJss8JiTPAzoLBFuB1qSjz2jwaSzIL3F+oF
Uezn38Y6qUCafG5R46eJFH76QJ99OxUodHgbm7nl+D1v9Xkk83vKgXafEMIa4sD1ulr4w5Gz5Kya
ViBrD75Jg7NE/DILsXiNF5VA3e6u4Slm+HA+2e3XS6UrTSV+ywGA3/iSgm4V1ZlUL8tK9VQXNQr1
rmUHGCj9Nfvk5wwKtMExr+RmEfoKT4VO/XIgmiQoh+Hkv02ibNb0x4fZnRJzSCrYMroWn8nq7snk
04HQUbTaROFV4DToeV1gxWXH1atp8Mx2iRz+5xJnGSo4FJtJr6myp3iIpXiDJvqWz97kx6TySgDm
mHaUCmXSnqGQyVuXyv6LINIznbHmkftHnpuEc0LNOVhVtd4sTiT+7TGCLTyW6AalsfBU7n5hcMv5
m0hjL+j7kkz3iXc2su7dEKy+QaRvbU7lPjFFHBCuv+fmYRMUWgJPY6B9c3jjeyT2KbOdgNEG9yAt
0lpq/uFDSVskBP/aNrsUsmy4W+p5LOdWb/60K3MFKbUCGGFQ+NjR9A/0UGWiDqVmtrZXvG7KbxIQ
GJurf/HE6OI4csW6mjsmCIZnw5P1/i8fbtPI97ule5WugIL3L1vzUiPJPloMXAU+i8qKln8GZKGi
nH2VBFgaD2pM989J/kySjc+g1EqGOFeD+c0eqOsCgBis4tBaSwbNo8ogeBvVMoFF5vlCh+2+76D5
WUvH5WUO+i+2s1NsimrB7UIZnOQ2Ml60YZtgRV+f/Dfje6VlhAVO/jTQOLxt/48bpDe9Xh6+HiCz
UIIO1tdgxiP7/EUNn4B4fHcNdBQwPib1/68KfF4VIxOwSburHLrrfnLCOD/c3C0zHiJ1k7J19HEE
vrFdS9UHvTd/lhfAyWhRTEWl+/EZaV4fQDFd6YQCfEKPXxS92As+MAQP4YSY9UDxJMkvf8cmmDwq
uMsEak6maYAsj4O7d7q8Ib/Jd90pjRVEsixAeK4ft0SInxpJWcR4+SKfgTG41O7gTDtLb6lS4Vjm
Gfqbw0PEIMaLokC1Hyetw7ttJT88lxyQBBAHMQlRqfVMz8nnIgpkDyOF/6GrgO0+tSQRpq0Jk2kO
Dtc9NH9+JSkFxYBJFBI7yuQY/UfSZPKRYQE6/gHxu6ps1oFkIilOKtdtsKKJ4Xv/njRVODQuRLBI
OKBkbzQL29wVvBJMahTnZcz7u6p1Kfun+7BXbpmmEEKOKggKPOnRdXuz5UHZT44vAWJGtdi6mcoK
R8idjdmcUX5KlxIMv3UIHLN4L7RpmLJHPI95kUPVFMyTX+QWZqEVFWbiQn1l4U6yqsFhUHBFE/O4
OhixiJFrjJDdq7WthZlN6GRqVXX7C/K4qHYkRW9/hLeaaew+x6vNAL/0f86L0R+U5UfUecPqcnzM
C1cSFdAXEynXV3yyVovxOB0lVxDBe7dszcwFPFMU8RpuHagBTQFqyhbi+wjvWSDdnA//Dw+MHJkn
SX4Vj+WRJ/EcdNjHnBMCJHJPJqu0tsf0x7lCT8als1KoTInHJj3ikrB+3ankBy7Do17Iw4iT7xkl
+Fvi7me55S5oH5tZaWRUzAp4lwea7kMUeN4VkcP89EupXmfpKrp5f5KD4viYkY+1Eaen9I8Ogyiq
6Vyv855qBk6ukO8ra5cUtcaaSqAOVqSvXzAHbfCyDSn9kNpzeuzLb95HTBJDzfHWETeicPw0hfq8
C1Ak66hGqiveZjENAJnfEIhHeT7OL6jmtokZb+A7BlqwfkCHGD6RuGSPqnESdf1JV35ar8IgfNIE
uCa8SjGOYPSxBlNkWlSa0OkaoKTeq51LNLZjM81OJja04DMG49Tl3jaQEQglgSJrQ5sf3wJ8Asza
A5QHp809PClIu0iqc6rKExZZYIEjwEkUuPD6ZobjAgVDlOjslDbWESlalU40uAsYuuBn0hXkzOKy
7hxHpeS+uK6u3nPgA9xoNoyA0EQWuRVCOkAeK7gv4QORA3/wTRMie0RvVfy7ZYCt/EQriEDnU04B
IiYeSqyX6ywLAmFIdVFbCQusM7SQgC/4CDmTOgRP786jEqdHj1OwuTqRbK+hMeeGXcpz6278wOcS
xrppPmifm2pxZhk3R6IO/xt09jmGFZKzzkljIYkd0OtSp3yn4INnEPuHAYq1ef/b50o0jFEIiV0G
gOMIcsxI/PGGdX9UupLetIlD4VoGWK1ZvCYFc+clIX/0J/n9XGmJmSxSR92htdNai0jHv5yHZJ4E
ljLSUNexMkhIyX3tWPH9cObQeFZ1rm3p1PeTH5UgmxEut2Rf54/BCmtKeoeWTo1wKw6fJVPJuNrj
V0yvYbQsJg+bWEDpbzc/nnsy8J1Us62+TdK/P+UZWi5gElSeaQBl50mZaVMf33Qjv6yfYCUW6m2A
0Ye0Xm4Qe7anDLdJo8FDCoNbXHbU5uyLiAiZts2scUK6ow+Cfr5iaUqp8U82dkji9tG2Bt3bDuvf
Aap12sD+4S0Pb3thCtBjU7ZTKDbTc5/tZUHHA9o67wiY0QhZvMhnmHxbort2RYr0JSM19IajKlb6
NamzyL+/Q5cNAW0llfZMnGVJOm7MfZIvFx7CLZyKzWgLC5zIhhMacWwr1VJrxL9/RZV8em8vcKRe
opY4Rr1+0fMcbqylhpy+2VfHuGo8oYb+9kL1JGGWAV9GBHFplLlqHQtG3F+RCanfq5cArh9AL7NL
eh0Z1BWgWu5l8CS1R+xY0i5aNBiBH+9sz9TkXQtoFZVlKeB2n1AX/H22xNE1qyIjcU3WLIwFC9S1
8WLc7Y/D+/TwkGqXiQyKLy/4QY2NoE5dsexhRVz+N5w+fDdx9HfI+6314vmofgla8ZZX6gClfZTJ
UOtB2OxAsO2iFgzuYN2b5DMCLf0UqvHSw/RWoiJFUNWh6vxpi6+XnEh9yxGORcPI4ZOsBti9/7A8
vnSv6aypLK3n21nU0SO7jNscUwo6ufK+ygx8EcQcnkaKjG6kZPm2YHnGH7DzU90e1jfWbt0MPFnw
odSLXMrxOaTPvcWrr6NOSYuC9MgHC3uy1UpgaBlC2BPfjkBH+uj6XU4GfhbykO72pv3kCO1V/Mbu
i0e0A3YhrhFj5meM9xRmWugmyZmd2JkJJih3wrY5WHjJLyINncCX2L6pZUZwP97VNHREC4+nrSpL
9Hzur+RXCpCY4vOmSpA7V5/uhK1lK31FvpLdGWja/wWlno1Dr080nAc1HWu4PNx2Ie2lQHanu2fB
xt9W+O1xm41GRgmha62qLhSVOjQn6Toh+XpFTlZsKL4mXlA+vNXV7DnGtntbiQ9Cm7uzduBVusf9
pIjXk1G7+WqC04O+OsSFt3HG5ltsyGxkb/wDYXaAdwB/V8lHP8oxKAG6q4CLG4CMrqoCYls2ESSJ
wmVHxv2vUZyhvrzxXcFhuGYCwiFqHr+2X67FShVGZw4yCq/XKNMQZ7zhraJYyFizEoZ8XTQ9ITVM
YxmDEn6wMUqcjQUowK4wbNL1fdu8CeM+zYkE0Xd/7d0TSAI/WjkkdswuYVbux1tpvxoymOxrLOJM
AU/AqsgtK1rmAo5dyMcHhRV8vkMrf4Y3uD21tJiyxuCGHECq4xz3ZSuvSlO5cI5yFZoAkXQNJHKG
U0pA5W4GCSRlQzTM4GjNflquFlJ9iaP7QxURd9WKIMSrkfNCGrHTLvWrLpPFhItgaOZ5vrRDLD+D
5o7X2cJC23S9iNnjuYSy0hpHrfsgcQOOo9OrVaiEUhpvFu7aKKZNcyMcXmmABBGMKfP8z+kTD2xr
sLoW8C4Mh15VWOG8oQ+fbMqQU1nKrbTtN1lKVx+qG9acEPhsPpmd5A6l0YJhKX/TjQmunXFTjmVk
Y4dMewuDXro6PhtvvNoZKhPGybGauvGMrQ8aYcg5apE44n+W/YhOIIsOqrzyriqaUGwJjZNC+x1y
f1Z/C71OSfI9EJld/S/dRFYJD+O8lWEgxnIqSFr0zQ8SD08sSzqYPVRERxX3RTj219vhffkKqyQA
5EQsrW6sIeVSYACM1V/ds/gKV5iIRwcQSgtyuus/GNXI0BVhQM72dmJKFYVlbz6X1D8ZvPBKWMqa
Na1aS236E7FFSqg0/m6ju7S2bgTj0n6MWH8V+vxHoKMZ/yL/8Q9Z3xKx3M3a0S/nw8zUGf7+b3c0
U8oaArj0LOI1a6dj+cWX26B7oV+u+yWZ5u1XU6LP+HTPi6HdYKI9RjnoC6P+J//QS2XwramexyZK
Qh5J3AltN9A5aEMG8wBEATA8oT0AwD9t1nv0SAjy+11OP8JmBvIB+wQ4fbVo6aqCrJqH+QYtBGs9
Jeyyl1phj6xHXh67i6z14OxU389s14Jhveql9dk4MiMLnlqP36sgyMPJ0MJCE9thAtkTPHatQXXE
RNbuILqdMRMhDTf/tnnbLLQ2p/PdeQF+YjRJ39nGSnsSmNuitSm6A/CsicriUFzRV6LlDmW6i2bc
6LIuqTNeRlvnUQCgUNayYAtpulMOVoC4SzP42jqAATyV2mXEh6oCiviuo+YNEgvhRNIXJ7UFe2ef
0bqQHFZNVtWbg3aT1JkR3ENrdD6KEpofvIuqVTs1Vvui/k3x7syeu/zqtmhJqMPENDvGnQa++xwH
IUtiQ6b9ixmN8v2XPstCp8+913JPcmoGsLZfVMuh0fiEMCrXqoPy354gO4AELRVHoBJTykt+Q4us
J5V0r0RoHL5mHplzcM+shoBsLxbduoucB96oyH6hZ/wyKJmfmcdN2HKuXXh0kXlb3E9FuAEEBXDd
cCNdFz/dgeAy45AnwjmHOPYkyI3O9c7xWK+T7rpN4/z+Ikpgpin1nMiqaGZi3Qwu67aj7EF3nwpW
RyzOt+Ysz3ADiKZAFrDC7xQHQfBqlcW2qKOwT5WoPkA/Gka+p7V75AaEUOfGx+kTFM5sI6h9LTGC
aiXMyn4XLYx9QciAwG1PH8wWVO4i1SQhQrC97rDbE/wooX2pv4vgq2Kyu7g1DsoR+5en3XXQXWHf
YUltOCAsoIPqhqrqGmkTsjLlpjJ7kBM84U129GukYlFrW9igQpDE1BB1jrOQm9s8bVwjHzOq9xog
YZMAaHzc0sDPIZehAAA4LWjex9Hs3vwU8SenXSSbVsiT4IjTTF9Leqe84oEOS89JAgNjtu3XK9/M
FuLwq8gRucPJZhic7rQTatAhkS0eK05InLDbG/VOYC2JblpvViap5fRbO174nemc5IhVqrSAm0XH
yHExCpk1Hm9HD+qUqADepXDh4K2nuKQ29mAbV5mGJ5g8XArwR2MYXqgloxiWhajFIRJP/7VbVQfp
GnL8Js9BSpcp358iLCy9gTmzuHWS2CZVy5mfNa4CD98cUAC+Lshw4zj/6nquubXtBHwQfiXVI2hW
DCib/QRdy3Tux3HzJN2+L3+oIYoSCPNiQwg01CJ0BV5c5k075ej1dBRkb9lpCirRBBkfao2nWrqD
ddNFnmZfHaHZujnjY40Blau/yT3GYlrSwC2RPz/MNvQhQfEGgeSBL/xdXlhG0dBy4ZkJshImvvS0
GReU06aGcRK98mJkzCy8CajFzl/XY2GjXTJx5H1weAb/eK0fjimCZrY25sH3n3BjCdVirsXVHaO4
s/yfZ+bazVIa+WZNYSvbqoVi1TlkNvaTRd9qEaPLvtxXMRC1tp1jDMRi/A8p4s7xmw/OebPGahVH
AxhOHCUcwphSmZ90JX6X6o+RIulSxmkKvQpgExRPPZpG/BZEc0rsdbvmZUEihQsIY2rqQU1UwOFk
iGM8ckMkmsD50yT7rnGZi+1upzTKfkYiO+mifAjZiczlDaiKENWxmTaPK4kbb+fY64n09Clmzxb4
ToldDYVwbTyuFe8zQ5kDta5VIU3vp3W986nJ82pmq8VvYOnW2WeC++4p3KVZ0RMYb1EgcpNgePpd
qWFpNeHt5GzuPnVoYIs2h5PXPUn7ssNrnGdjnak3I5Ov1xokd0Q/FxuWyUW+l2sJVIp5mZmmKJav
bkY2O5nq1PAKfsz7ankVIymzCxLZKeZv5MNp1ExAklbLpeHJBBErrXaBodODYV3O4dgxwPnx4ow9
RF7MZodhwvEp+Vtkylfc/tW9kcuHwkvxOGlJWTpJaAkPdQHiSXxXpvndccbtQ5L9meiWUpKMPgdb
YUSj7tRADyXd8tqoi2gz72kiWsjD7Qx3lRakOEpXfn/o5BrC2V7CysHxstdj8eWqCoVDsMH70Fh5
EKF70TjWZcItscfcGUk9dqD7ky95eV3tqv2+/Iy0QtVJDjTwQI6rj94BZRDQQ+XYgqq5w8BYl+Jo
dbLGc+KsNgHGw3BAXK9J+GbKNCcI8uTwh+3U7icy8+eHpLoWG2N24aurfblARop5gsnaX68H5QwR
31SqtVBVDfHD2Mlcx2ilX0/t2RPG7dM0lMKY9gOViZuU/KFXH+t7zg3uiGKv4IkdarF4HSd7dQ/i
BLoTFaMresqpLFM1IPJl5zCioaw/JYxSU5XWQMdqK7NuSOLX+1asuk5nBSn6nZrOMnwol9fGQ3MC
WJlTKcBl1YPIqCQfS+mxeMcw6qSJ9Uz+UdB1t1LIeNjTFX0+EtgZ9R5aKd/GfzWq23iLWQHYTJPy
Em+XAYDeeS8e0EnpfYk0UMQA9yKxX8iYigYD1VSW48JSXY8ZG01HAhlM05eAyqZ4sUAjJ+5GNTlF
uaDOMxmHQQ+hKQP8KjfK3zRHX6dzTULx7Bq+JuwDH8tc5JP8bMYcJgxcGbxegDK76J2+DVdonwuy
JaEHlTO37HsaWqGbFlQ8WaA6FLGcY9f3PbreRdQTpOKBKjk4mdFHCIM8TizpUOThPPq6cqhtv9Va
0EGQS/JEAFxiDt40JK/vyu2DXsipylTxD6dhv0kRJAiTJnmkr441L+vKAp3fg0OZWTorDml2OPdg
WmKhENmPWOGwbsFuxRiRhy9ZJX6SdT/xnoW5GMPE98aAsWuQDv3pTV8fp+EnCF69quHziAk0EUnl
Bl7ehpWeDnSyUGrxBbEN0/GwY40cmWtj5m6Wr5lFZgXmAlDwEFjVGC2TyH8/Mu1coQXdvjZoUbIO
iX0IVt4cYGt0r7ygILNzuCqvxmUtKK8saMKHnIigeaWkkPs0pc+dvv4AA80mIrYjqSG+wAcOvwot
MaZla02EIpxSaK5wkJ9igA8DguUm92oUj7Yn1jtDPV3ZP3iReknAcyI/Yweqvn6IuRZaTAZSXd87
1aVemMy6h9gLqYUjC0UHEsUUqnxkwS1/ZHDnb5CClPmnoIryVveSOsoGCzoZwuxpiiS9rUat0aqO
e128UwJeg1A6VhWqMzIyJKQ9Y9vGW4iXnI++l55Oq8fH+1HOC0XrXPvdZBs59aK5Mh3AGhRZBMNp
NXsQbP5zG42c1YWIkzCMXg/yqOBP30uLVLQqsVhw5IaiXUaIQJC4AGnvOxpHzQsQZZ++0iBSnuyb
M/O8HDwJdXL+fueK4TCykX3hzKISrOVYT2fpY9MIDnh6dBf1G/SJyGE+7+T3qP4umP+M2FI8R5ec
1yAmpk3ksPMSEn8oWQ8fMVJ3zKS5emWtWvAJy91lFBQrvG3wkyhQmAeZOhQV7sjGIJccSH16M61a
ktPrn5SISZUcI2D8c4wjwINOH3cm3lD8uPz6cPyjVzihq9ctIsOoidoTh+mmVjP1F1rdIJkAZmOz
4qKy1IzcFdeXkK18A7uvZg49AugPJZtOivCJvMng4cF5NEZuT9Wy+kAq1Ju/1UIrKaR9nF5tjiE/
4hgbbkoX4T4PEjzJF5XOvhaqyj8yvpv2dwbLYhD71Fm8BZH5Y+A+dDcDyLWaODM9kpNdMWn5wgeI
0UEAZTRB85+Zm+V7LhnyBdL3+hObWQAM8Z3FKk9gyKHR8K28GVRdf7kQHtbO/+RSpaVrNvNsR8ra
01cU1Tvg22D3Ebt5fBHb5WikLhqOSj7MfNK7BflR2QJ6Uc/kwefOqwh+8+5mW5PGSttCFF5w6/6/
C5idrXMi9GjvLUiqsYaonEyQiAzqEfAWFntjIgXxnrVTUFYxp6zWdGsC1JoxFPEVyknNishVhn/x
435YnXix8QCMeuaxqwCLYnssQfzBzOKh72yZKJKqJZkwcdHe2kmA2xhnCJb+OwKi5rhPPaK9Ilcs
y8zmgz8wnqI2stjMa6XTxJaI2Sb9leAdCs3YzPdO33tfrwM8Qrc+IdZyNBNXHpb4HNwY5KEkJh1d
i9ziS6GvHCalOqFAG+uq4L+tImnLr7VSKuxSJDzdsGh84ZUSN4yomtxfdhMZ6VDPKeb4yVaNFktc
XgSqZUnKSeEzwWryKjg5hVdiheDoW2gN0b5Pe+bpTnYbbjG7G3cwPeCc73h4YMljpoR/43UY0B4E
UUROWizjt5OnHrqYqCQzRXPrkU7pdR3p793n42N4mtXTvJ/T/bJHW0Xyo0Mr2uF3hsT9PQasBO3P
RyPyrE4hEWYVpydXReS4jUbgLRtcFAAwzahKb61em0REIqF3P1VPhJAOhgS6ZRhOyT+zDWPGTIkC
cPDA6RzaIEk3Q7L62Y3foeeTfRUSolc/tCCRQi6PqiKJz2MiNQBCanNAbqWDGKS5f6PnJhcvpFrH
/sHqZwj03YZn4E9U4G6aBqhtxgqI2qxoDfl6DPf8ysQrCAoIoJ+hrt0J83+jLggkytdg3gyyxHpS
IsKSWYqiFqFIqps6JjzKfRwAHvxMyXqsyPVFVQRiWjRMiPm4Yweyzr303cJCglUR9pjy/ILubvip
Vu+Q/aTwyLPIB3xUwz8t+nHhj4QuFx/rH7LbMibXBKi0s48A8wlcAe23hyhX3NebZi5kHtS/YTFu
WPvW6RBAn/uTqC3X2oWfJVB2CARILjfjXd9KRo60W7B6GGRsXTzMHQF1031nfEIZx3gyrZy6e8/U
ZUgLWuNzsk7PcPnIx49XMcPsdZJkOqrB1tuM/dMctKhBG2xMbd7Jk2GYWsiHL/PI0K1GGPBhZlNq
qP+77tEYUNSTlYjDR1ILJxHf/RFB7lS2CADxHqP2SJw5EhoRY5sDB6qESee4YIX4alZjQh3tlTZ4
k3zLSxyvIfRbe5yZvJx+WzU51a/jlThtkJyigJayJWqV54z8iwu3URS8ggs0cNJiI/sPzNU2t6bb
o0Sim9In8h+8Gb4kKcKCHvZFewakbPTwe4eZWEdnLoxM+650cIuO1heKDaFdUFtVQDt62viwZTc+
RpbgWBE1WqMfDdsFO1TcyJqT+S0mRMVp5YHPgFKEgimqcUxWMFTxw/bb0Pr55eIYgPLCtMZmFmhz
gutu4Xer9LmFXbJkMP2teDH0OhNFYoeLRWhoScvTSRUXH6o4iuhh8COQ9mJocdaU5vbfn0rkxcL4
6BX2T+vc8eanMs3t+18j16jzctAWysug/AhGSSBZBcjFltDmqVdLdHE9v1hspgAVzPyRe1drXhJa
B/ipeshPRV/8i6qd9fV/dmP+n9+5O1uwKT6+KQ/iz7GX+X8sHMQo8KopKFTTgwGq0CM44HAVIwo4
YieODw++Qtb0wl8WxZ7yZVXR/6Rpd58St2SBZ5AOg+J2eIKzZOKSzVWxiPIh3Psh0DkySM5Yhd2V
h8CRNYj0zfcQ8W7L9f9m81AgBngJG/PgQ1XgUu6vJ51usM6Ig3DkzOVpU5QDL3DiWXZk5Hc1EhCb
DrSFA9jd+DieS7R1mUfB4PFwodHnE87wXOptwNB0vdrmB/Gr0P+GOwq3l58gFoVrcLn4ROP5fTGD
N2TMextYIq8qQrLu4nfWRaxjSyHHj5zdy6twoFork+3gjctyYB7g73T0Wzx/NGKEP1gZVikwpgWz
62yQeAVUFyu4yTUER7eeFlAyu0jWnsYM/UZ6WwJaXi3zv87H0ojRQWRxHDVSvl5SG7lHRZtCsjTX
7Hldv/r7A3JKsT/EAzVS6R7h6azHhO0eKzBoCKPWap0cZVooHgtvCIPYHqGK+QfSrqNsLqA3DzQ6
EtmHS7L7HKUqGL1ax7/kAmnQBdcL4TWYALEByz+pgfApOdY2ABDPM/VDmeM4xhlmkd4ILzgMRY6x
JS57Z1KJB9vuCela8Oi8Ye8DjIaOnR+G9DesXtuzP86847eUeeJHaRQY0sQY44rt539uMWDjcSNd
j1JIf+2F9wzkUii5rivD5Cfmw8pG/A/xtDEo8qy9TBsjz9od5+wDu8ClpsPXNtqtIM35wVy7kqCh
MrPsJ8WnedCR7Hk4phUIjephnCkeBDZx42YPT43v3do5rsMUlrFB80fG9efyjMbj8NlBi8TXx5Yw
g/oZWO9YSKN/4OFcZ4Ss+TpxG8aMYAYSl6AaZmuboS0W8IZuDPkF+s/QLEAQADqQYg93ZFUFv+eo
gQmEJjFPnHloPY29d9Y8qUULjqreU6Vuk4eB0RO+yTlmrzQeR0E+QtaQ675xRnBcz+Ou7hs/fLX1
K6nWm8lUcgG9Wj1KLKoiyVOvTML2YORqH1F63M872OaMVBmKnM/2yzPbEsQNa3tDwF7jDGp3GZhx
D8i2s+/MahFbgPiSjjkz7FokbknTOhxN4j9AlBRTkheorFF9UQi1gdn04+Er2JAe0tVKoUgrqc58
npKtqZ0BufJmeQZpEfZAwoERA10ARS6JMfgE/CcG9zRZ2TBCuWyQ3UhKwjd3qb+ETCTIZcb6uj3U
qvgSX1i2GWQgNqKvBLrNy+C90ALcCoBh7xsTVZgtM8QjBt0eg/i6b6crIocK2h7I8zdRJcFB+xfA
/TyiYcsyUjseYtc07agOgjImbU/Jwpn8oGb/hmDKc3pyi33iAGHAasMUqVAzF0hH9PQifHQsDsDu
OL73kAMrd2TvgWbqOzU8qo+veAqtmmshtChcEveB9beuFuSsf6+nR/3GE1dOe189bcjauuyAF4HY
WMAyudtDAoiUT5oTkWhusIesU0x8Xi4QB96qyHD6qZIYY5yQ7OhsFU/35lG4BBrUVJ+vDTfvnjhf
5MqMGY3ohRWkV9XPTt1UbPLr5vvtmon/O4NQge95NXxLe8C76oQFN+A82jAekhzFhSDK3c0/An1T
Ac4wLs62TzN4DJHU5KX1JFMisXeMIlJZRt11XYYOTm7qGLkyRPQejv7IbhL8XSy6HmIvHerJo4M6
RoJCghaePyeHmCt9MWl+UZ8tOZzBIL9HDoz74OcAuCCOUx7zLfJ8GlNHlTKZxukAsTI6MHV/XcHU
dTvcI7ssLwp7n4W78V9U0u68eFzsTEn/EjZy/a+8m2z5ywGDe9E+9hcrTlCEAvw0RAZ6NOwuNkKc
DUSIKoSOit4w5+K6/SG6nHu/wwFRF6rU0E7x9eqqdfo2BYdYK+gcIF1s4HXENKINSmK8N0uKHaPH
3NlMEzVyXU9FhNPm+DZD/Nl2OlOZdli/NmFi2RAg+5w6AJ09jZu6BhLdRir4/uss0OfpuSxvFt24
YICR1/APHepIdvuhdCnk7BB3TTLS9TgyVjshB5/JWH83JAFJ3b8fB/j5fgtp2ArtOSKD3CWketQs
Ot5lmsw1jxOJEbT8EmozoCi1NlXreGtFrkVXX4GFFo6sXP3qWD2BTVHMBLQJ9Ea6KWJkynYVVkim
3ucMxIY03QlXHLjV/RqFVgb+AUtBaZuQP5aB218bAWokcI210pZkHyVc1OamYqpdr7G2y9oA8CtE
f6AAao13WIz4evz8F6mwL67WwuS66mch/MTC08IHGtX1PJ/hogqsCtb/TTDmNPID1faVHrYEbBt6
kn/Tjq621Na3WwuS1uqD/AJQt3gR974OW1r0fLSDufMlxBiMauFOD0GLCjmS1vVdKDIg7qeQkay/
RhNhKPAnGI/VQdjjoSDTGDTBZY8W1WZfw/XsXLkqYRfSxlzI9aiUJXe+GaFddB/FWkp16YAfyOYg
lk/As7cD+MpMWGgeZxMn0Wu0WtioFiuRYdaJsQIt4rW1RRofiZo7Hvj5IrHATOOqlzxaL50sj/d0
7XGXGU3+UHz/T9XCaiRU8oXu3X2QbYH7FpY44CMe2+k6+TMdcIRrje7vpt49pUbnOHuNDpRsM9iW
WV3xxVXeaLGMNDlU8ZxcX34jDpVWRNRVDFeem71QX0DPdtkq7/Fg2NUbMDjiwqBIRa1V70vfk4Be
StVm6KkiegkXaiHNfdrTdfXiK0EIPmzCHz7fRN3DhmErmOyXwBl1pnMJoRsNlhgARrb77LXqxzlo
7qcepVpICdorxFVFulV6IWtkPSwlmzv4TGN5Mn+QAZtkFlbbkgO0d5SaaxRwJ7v4a0oE4Txqpk3g
v/ePeARrQGuXnXM05E+zuYEO07LQPjZ5qwlwY68zEo6gAfoXo7jVw9U+XpucbMNw7ksAaG6hd8yz
3v4uyMc7z6lEFFa+g5XLC0EO7PSeGcWzaFWANsG7CtK3/A++CFUHPxi0L7j2vRjZGE8032MNJZJA
SsPJvYTkXDvEwI9o0oe2FKuRHn1kuuWRx7CxNsx+5bXBrXAIXNTGUJ5AY67xO+NJ9WK0VwPlyjb6
wMyhRVaYpo209/OU+oXXh/G9SirkOKXjFd8pDH2Jj+tBCYcc2MzWbdUYq3YA/MtXQ3UUBz0n4E+P
wnreQoLQwcwajXy7ZTM7M87PKjGfc9LK/s3CtyuYX30GXrkX2ZOBArpSr4IEj+7CdYohPA17qWjV
Skd1YbrMbE9mNc4xUvWx/2DgOl8D2ADxABcUmV5wS2oEcM05Ktx0/FzLANK6ekFNjhRRXTc7ylKo
ZwwTelOenpnMTnAvvbG1b0eGeKogpzBVHV1CgT6HhmsSqEtXFGrXb1+7/DMTo2SMzDUZ6YXhchf/
wHJHiS8CwJaJgZIGIAtkiAOjfA0MCHXdJbKwZjFqv3In2TZ+oZuEFfLCd3I/LQnUhjObQ9bPaiq+
FkQVME6MyjqDrSN8TtRzRRlCc5xH9Tnw/RoOOmvo3aROA1SYZTZCr8TgAazxVCR8yqifSxdCng3e
JhOa2RHhlWFwuTRe6tZT/UqAhefG5LEi5EkuooqWK/kedGF3SCmS83vtSvGDB82aTigC+WjpjBi0
5+fjIKxgg85es04vEbkbIWXrlNE+KbQojvv83R058ZHbvRZdJ/7+J39B1V+qrwRst36k+EbFP08f
6I0oLxL5zNSAQGh9D2ZxqaymRMyd6/AIrTyrayVRGZFpYb/XLt7Q/CxXkO9/ZZKwFuypdjgp2GsY
cPbL+KTRPc3NwJHPawLUdndoVgbMkj45BlusRfrwZ5JHLG3sxIMxilLn4wE1+a4iSyn0VfAp5OvH
pOOkXdfrsnEyFyZJetYes8TjdsWUJF2zbgX3DYdARz1ZoCXH9TCfxI27zojIeMyTDq0KC4+lDmwD
HrzI3/MB7vuNUXsBKYmMoxNr+eeN8SckVgW0Z0aiPj6RungB/bESeX6FewYUzvWrzyAVzL2PTugh
gl0DIJogjoOiB5cigdBwo51pKaXkUJYAnfBFKIDDlppd+lsIVFf3MERxUDLG7JPjT/2AkhpwxpH+
Ffu7gUyZwaQD3ksQNNuU5b2Gb3e0T5koe7LmR7Y3GExnCISSd2YTCZ4JS2IZhwa8zExgDYLGQFq1
MP63dwzkaj0U0Pu6FF4sGPcwshrZfSwen6kPcU0WB7fPkqqtfNPA5r7BjqA11b/3K0ebewtB+9Ge
nGiXIEH9enqWsdXXTL6tRshyU3HkX250EBzaRyCZSCTEVJQMm2wDf0wp2LAG5ER2e4jUk0ocPu6x
ZMA+HGi+/Po4LgBSb7yYqZDts21W1GgEY3Q2HsR4Oe3uTRUDPNlFsBfOgbkLkiX9LReD0Y8n+Rlv
6YtSVyjaq2/bDW0kkQpFJfyoKB9kMcL1wtjvoiCCJcsh23fPXxtVpurb8F8RFIbdG/8d6yx0S8S/
nX0YGzLMt8sXnZ5PpAmJAAqpYgGOwevpnAs1Ghz75OOUNNGZiXgii/hT9G0El2Idg6PU71CK77Hl
Dl2vKo9vcWQQDjgWj8w569fC7XangKK2KGQSQWHKNkuoSHqzdBE1og/Q4IhUU1M3g+Pulg+xQTfb
zO970pLS8rXP3/WD1g4B2adKH3PcutN5aRBBfy3ZJauD+lU9aiaABSS9JtQcCh8YpeQ56JaShQId
VrP73bOptrBzosFfCFKi+cOFlLIrDtmHNNBdQO7LlXU5idxRVQLeQ7W8rhqOIu5gd3iR19JoOUgW
UPvPGo9B56y3x7Sh3re0mtgP7LFHvv6IMm9wKe5MB6YTfcHfNhvkLng5IX/BwMM4pmzqfXQduvM+
egvJJg161c8VKjI62+gedLslEnU2RvzNx3ZvXMfra/yaK5Y/si8ZinGNLL8hvhUhHPvjaJ2Ve6Hk
hDjbOSjoR8hHvLWyVNYcQYfbM6L1ctriQ1D+BgUNlO+SCB5P64PUq5cykk32E0dQjueutz7XZ+sU
zXq0oRsFaCcdWs3mHJ1FcINw46voCMp3yLQdhyUXsFWyBCTgncLH0cDyAJ3jrFCUmN1CJRV1HZIk
frGdApQNR/xT3tO5/4+ZDYGyxi9AS5Dt2Lih6REMdgXEvGpgCh1DHz1pliSEBpoheyvUqsR4ArbM
Ob/2c3TOgJkVYNcCaNOAYNaDvWoYcTOm07iz0YVhJCcaJEa0XNxR3TvkmHr4sppw8eRhNeqtRznP
3z+WfFxRdL/ovftr33cCBkBvISbVtUW24cgTBQB0kLYrNb8KrnX88g53VEKUCYhG6w6SasAgzTIW
BR6FgJW8RXYTd/EdgHqQ+1NaBjd3YFq3ogma+H6Fb0NtfAoZNUSNr1iForQjQU1jCOGWAlnwpmfC
dgzFCFWqM45b2Hfq/91gKJa0uvWY3phc18z61zwbFX6gYbebGa7DGv2olVV9ILrJoPJ1viNDEfeV
qAsErX/G+S8gmhvw+1YEPDAUEP3p2S9xykQEe6ETfstrY5ebX2cQG1hebpRMQhsLhpsLAfNeA625
rdaqZQ/Iqe2vU4ihALC8OijFaTIfVnqtTAD3G7Copfy9ktiy8JyUpBjZrEFYhooACKE/JF/EHN7e
R3Xkpce3/Ryw5BAqpZ2cxV3sIFB1vBPKTuaWolqj6lfqU31eliLu8WvlDl5nW9Ve5UilecHnnUSi
4tePOsmI6d0Nzu0XMDGGT1QZ1vnS0jF3eEn4EH2BvWr85JqRyGGpOfz8DepSW5asuCSwf2OP7xiI
autk/Wha3hKmWF4md2iL+Bf2HYRpakyuit8ENTYhgmd8i9hLA+AB8JlbLzalVo0iBi1SJvRdBU+a
/0DNBzd89oMq2OGb6THhfSXPM0aAN+Iq9vyBqeJqnNXuJ/zSQ4lEey1Q5/AjJ1iE1pYJZ5+tEAEc
FwcQI3aGMiQBHizG4TFy/AfKbaPgdZRCDNgF2DpINOjHvwOIf8uR7RGxbw8+fzezslQN1NDhsF9K
eZxxsP3BXRQAq33kMERErZ2uzHcMwoDeuJ+wg9dDVWpfSpq3qRswPLLdkD2/MqbS5q441O42Dp3o
jrxJaFsmhfecTwJADi0bEt0drn+TqnVDVtERKaOFPYR0znfjpK6SLEwtNuBKbwzedymsmCJomKJR
Cxkq9lHyaLwFNKn8jdX+kXEm0RyNyKtbRQNqkY6k5/5f41EKnOohMGqxVOle7klkEU/gWA5lfV92
JjS2JE8GhwRcqYRGsQfpqcg8rFlHXSXXDm3mp9K0QxBNtleoDtjCtX2c0bo6ShsJnxWfYU8OR6Et
xZWl88GXPzMri1NO0z+pzdZmSz2NGXTS42/JcvlQ6qpxqJcN4KiDpqUYPyvCcBsvLkaWdYfOhV0N
AYHqSH+kDmLDRGvDqalsgXs2/p2Q5xvln6+X/rdA2X50mUd+VwYate9aogdaIyB4QkKI0MbL3FVm
qd1sfBJiDlegYNKqLcSLITrAZW19Mi4Ln7nrZTTtKbjLQgDDLsPchYRvHVp93C4TNWZdkSvtWnYN
zVI+7exH/R6yrIb8ZdDqP7Y+RF8IjUjokPsOVpuD2vokE9GhQTs4xnQ/c+TpB5+2gZWHUzRAB30u
3xCFvuQAZQKczPkucpLjIGJ8mmO+GCIh5qSV130qlKgbZHBHxFC72hEOUnCJK6RbP2MQBrw7ZS/M
OAb/q58FpZUA/L9BJ6dxbUrbZT7gF/iLp+Ix2tmgL7h/g86B49VEWK5P71DzRYDbA8rFM9v2PFMr
ZMJekT8o4Km1hOqqqLclbfycGVCILIkKh03TZ3t5a2ono2RkiCE+KiKYLat03FBPyf35FzzrGuIW
uE6Og6TGHShZhjh3VvUkAtNtuX2nqgXeHLoWBAa3zSYCHz0M26IhDuMF59of1pTj0lznMeBBmdEI
JeMmZfuBOXhGxfYK8WMT3Nu73d6HpoLj3mYpvkuqWUyApzfDzckPNTz5Wyk8wBfBOikwU151Xd72
b/XDKtEcQwm3vQGrmNlGr5c6lo0TskL5DsmAcfc3ToBydzPJIYR1LoskyfYwV8GWmTIWT87IHwln
E8L3v9RZXhLCFpQ0mSZwaF5CzEUV5DbNxwlI6KBeRLz/JyEg3/HAKghjyPXguon4xSRh/KJTXXr9
TZs3veWqxu65q8UrmHMYexwZVVyxYQwHKwPPUQ1rHPK7+DdWxIp/H0MZYJdNaBpoBg+Mt3OYkBDI
/Qh9rP6H3QFX4AQh8/4LzORu+Evju8HWBUwceXcOU2720W2iFSn2JiIKsFtGQb1md9o7uA9eQd0e
fKjOBjT0Krvc+UzvGk59yFKAU0vSp6sjrrEeupdrlCFpETMaO/5IcRgmGxY6D9SVpGSiNpdHo0fW
9e7uFE9OyRKjnQ9AzEmtwM3OCY8SE3HkbeKoNGMW2yy6iRJKqd98aOySktEaKt5cvR+7o7N1TR01
9S0ssJlNst+Pxrx2US1Ufa7uyQdrgI6MGkqrp6OhnhMgMQMSsoWiKETo+ENgYpoq+SjWSTsrU90k
546Ub7gfPRZ6rnCy58fKLkj/Di8WDoYLNt/xKFQEtM98FfodJg52QTa301lC9rb2D06xSMD0LTTE
34nrzkbbCvaKkcJ6uWBa9Df9UyXL/p0fbTdu0dfTpJLFZPq7RsquJJBoDNPF995WgfzEV159dDZb
xv5OksHlZOVHTf72LADkJ8NbZVzRLplWBsrWEdIiq+UGZ7ptVkQJezIOE0VWV2fiKnpc1a84ANFq
Pa/yJmG1RyFfiCQQdLZVZC5YW7r0eyF5gqQGCdyvlKaW3tC0I/RnmIOQZLikDgpQSgmRd7c5Py8F
6UyiUTP+HMp1OvWlG0js/8/w8BSEvNupcwPJboOQQuqwJgRPwlPl9NUmsd5SSom74E5BUPdwiNDR
6Ce9Wr2TvgwdQrZUzMinEWDbqKkD+dDNvgBtwY7FtQEC/AYlRn+aXYTsbrqQtmi6eXa7/szD+w+/
+edNQP2QE0KcGzlw+D6QG2g42A+s+xh7cjFwVfLEr4ZNvN0SAkQQSCdCSnTqoVtfz9svM428hMty
5BfhsErRQa4ccaJjz6CB2rME4BebiKpc+EIiDHpkmtwRb+CCdLearqbep5CMKMydqXxZxW2RwmQd
WbAuV7vAvhiJLqGKP23yc3OGlqjt5p6QdX2cPYoJhue2dn2Tl4coht4jfCza+1zTppeJ5JSg5XQn
mfSwopQPbFkeScSzkEZu1269VyioiDT4+8wnnWQyKBBUxDE8/cyHxDtuzIBcCfUVEF3ltsFRhZep
BNyX31DO0wnTc78OXJgrZQVGynkuOq6uD23rbSXtOSC7KNmt24KGbSQqMe/5iOgOmBj+yVlWHt3d
m4A43UErc78pxlgRstLNEyPp4luX7jal4UWXZIrQjiJVDxmbQauUV89KxI5La6F3nYdpToLG8jOc
tbP37fH0c98HszN/HHcGFisua0drUHbS2+uAP7elm+GQS/NfCUbcln1ZsKwrIKIENdeXQ59yioPg
bGUK7y9bdbGplv14sihLF4S2fOXZGcCnwRuouvovTCIz6oJmUdZIPEZ3Gf7CvtfuXDyPc9fkaj7g
Dz7HgzNlIZOfMtgtQ615MnEBVlZLfn2N/VF06k1qiBUB4INYVP/XTKJ78k8NPTEl51w9eI3TZGm5
NooOuAoaJghvvocILTkmX7Vs/G/i03X6GQ572c8wuKZrm9SWX+9Sri1sppzqEYFe+aT9sRb7Tnvr
CyUA5jaRe5uoX5QlDS8MsWj5DVKJP+WYDfMKGRS1taBk2bkpx5PcgOqAzhrCtjLJumRqtKLq37Zn
YKQ1VSYqREgFOhfAzQ74Uf41G1AJUx/SaOBhS9mXEFD/q/NNm84aKn+8yTBhxSCnA872Bokncniq
kYu71y8+c+B5xXkz5V5lOFxy8V9LpYfoWnTpQTUhv4pzEmkBUBhncoXv6XOx6ltvavlJpcGrlXwX
PnWlXnkt0mN2MbMC1uyv/bWNvruhHoi7OFFRVnaBVvH9ASTbJkkczfXPnYHCgsxeTKyRf5bWcb0O
pC8tWJgiqLSk/SDiHWIqntEByl78ZjHBOBlYmlByFNYZsHrKXN6pxAta/Tgn4CALW24PehsRQA9E
fXrJecZZaHYfKvplP4HUVwXX4ebtVyDwXgZWwkMQaCGbud7vOkvN0gSYe5af/F8irctQichdZnCA
rOs/OnA/ogh/6kyCbXCzstVnqbet7yCiOwfHRaBY9Yy+NmQYmau3F3OF5aK7+RsItgDu6jnknlMC
RLyIlintbeJDMtT+YXe0faVbmJgu52/EKDFZtUZ/CssfeRKGk04ucGdz96MGyR7wCc0GTcrk67Xy
oSl/T4tCxwXctuQdAAa8k+TrEsIjWYIPDF9DveJH25B3ltBd6B5S3fLf2/C5Igp/5XKZ6U5WTd3h
a51+QM7vEfkYRnRb0K2Qsl5dChRvUS/wRmX81wqKSO+B9Mot46ybFtoZRVJZqPnjhmEnTkWv076t
2SOwcNuQWKI2EWXCFx0ovL7sChpUAbrSBFZZm3UmC6rExutK18UpyrqDfratrpPg7szB6vfgJGKZ
AaNKgi5iXHF7YTR5CsQPvjabrDUOw2K4x1u7Gs5IfuUH2GMNk/Pib2vRcusdnWK+KpVnVBuOGWUf
3zFOONIo426m60lhJClbW5clSSi/21FxwNXTk5kgTZt4Yl+CpW/3h/D9ZxOi/MfKWDlprNCgC8gm
kZzMBnGoLS5FfIHo5D1eXBI4WkrB1Z2qtI2IHO5ww3tMWL/uW0dHooVpFx0Yu/tljRHz0yR1jVG9
OaWQqN9TJ75V8YUFfryVOmpGbJFOqjAi2FDAdnw1vmU5ewE4IHobZV8CLq1qxUMLq12nKQ9mntE7
Y9F350hdVY5dRSZHmkt5WTzdegA7luuCeWVKUg2t/qxWtNmtMylImyVqk5HOpViOmoC4bQxQjMHl
8SP2UcRhFvJBGXfUc+tTpKhRAygAHPk5Z/cvHEauVP/jKk72+YLg4Mhu7Llsfvonhq8djoy00q92
wVPpcNTK1qFg18Uoe0ua+P1Nzf0Y1HQ42HR/CKhBvxMe/LybHYGrteF7bMJlRM1w6XdOef2GMFh2
bzctC5dTn/XwKEiEiYF6NIREt9PvsFn1moBoBYbyz8JaFHTlxMOWjst6EsDw1LzQE1cxBiqTuy7+
amROQD1awhcN5ffKhqP95ai6lGcCIjIBAPiPIE2d4amcdAKQyRpz90Il+uBacxz7Cf7swx54puy2
FmrLxrPgd84qrkeCIVZy8yEo+qb8vH+NLt0pfdz/5v4bTaZWkHsXMpTbjWhi2pf4nhbfPgse5Uy6
l/JEzekOXlzB5XhjdUqm7lGcuRJNgEnGUbh65n1VBQoguXTzY2YDf15/YwNBFPGoBz1sIhKptMz/
DdhH7hBbSyxqKAJDFtTjBboeIG7EFdCTLoc3tc+DZdiu2Iu4JoBQiQDoK5HVI21pefDPvl/8bTG0
EdvM45iTvGS2RdN/z72bF7m/lWke0V5gkg2Y5uB0yWXI0qMwxPqrTk7JVLrHJ1zCGdjB1/epNWt8
dirdQuYrz/Wa2DoMX8r3BaIN2zonEchf4itlW+p6ychq7AL8O1pT6/0sinw5Q/+wWcND4bcZZ6qj
naIlaXviJHHFT72U4hf8OZd/e/r29fd4WQyw18r+DO1Zgh7NRTan9qtx5dSipoLizjR/sXNS6u1L
G7ZNafE12MBsJnmRD5l+wXQl8qteFGUY+0jzDbsO3jp0c6y3J3pVMYc8S9SgvkDsA0v51fRvRHd6
gxCtMdbm0YssQhH6hDPBizA4VxpBpW7SpZ+ipVcvMUBETdzDSpF8QAb/zV2dfKXXm8YcCptPc/4l
PZ2Twr3OMmJGRfk43HSqC+l4ByFMusi8oX0GB2ytlu/c3IPwLqhUqdEwUrKbIB88gSKswjVIglcM
5YeGgdogr9cBsKOp8BUuJ6WmAq/sPQ1bq6nUH+I26sW966exaXJoA8OU1/U2fVpOZJiXokwxv5fu
WQL+L/lKXv/F3P8awhL1dK3fhI9HNxFUE+JD3e4DrE1rQTO/Pd6RO+hQR/2Xg9I5AkGnZ1UTkZWR
7hXS3+HeWTD2mROz/qAjm3u52De60/yTaCh5reU6GWPshNBMXH6bZIdAi9X4u7StjmZEE7HP5+cn
V7GnNEgPMVm72mIcAOaIwXANptIUPbUHZW44ouyOPuHwyR+VjkVMOgGajVX+NBcT6/9ubmBH4OmQ
Aqnrk4SD4KQDu4Q1KLQoS7Y0VhDaHvfpd95QSfqegx55UJweeCUZT5jxyBZV8/8m/XORVeMqcXDw
3b6vsxRK2Lu4BNzlU541KIeh/RA15VxOodQK3VryOS1Sj2PgVTqspuUB+T2iU1M+QRWl1wiNjiHH
bpUwHutqLcFD4CuvD3mTPGCFDaUGlqBovweTydiMaIqHcSHiEQiSByq4hFuY4DuqhFbFq3yZZ3TL
9fBwfYX2790Djgr5lBnQ9FaSWjtho56zKlkIKjKCQP8wtHsxAhgjWSYPNkqQhpsMGmFoAj6UEfdc
5/AVS13cb5E3W3tbtN6tUwub6L00Rv37k4vJ7nAloYEht/GrijHaCY1mNfeFy9g6lTtS9DetO5kN
C/WAwr1pqHnoBMi9//ZLH1lGCO62cNZZu/TLVfr40lzBOWECpMPzvJ9WNvJHtAsgubj/vrxQBmh+
HrnFTR3m/Df5jnudwvriCpBwcUMWCVo/ExzWuOgHOW4oSFslqduujyVf5JByCXWd0lMAFgUc4/Sj
LGal1lH6ZY1pSeQwY285IQa35cXUHjkbYFu5OPO5lZWMLAtvyXBaLhT1L9osMwJujnOsMz323gYP
tHAkYvi8LLFHk47wcWp8lMSSQg9gt/AfgNtj10nuxkI2CcCEsdYZRHMuQiBp+CrqAX8Oi04MaVLw
pU/3UbCUYOgTW6nPwkhdyCmpZDMJrvb+Ncmp+XyYwRYB8XmDwAwVWEgrlmnCeg4lOcT0E9Z4tvEX
6IaihoecVIRlSX8dO0r09SXIT8CYSxw1PLNjutbHI9DxKu54RHun3W8pk2EM80qI+GsgEm6qUhH6
M7DUk2DlvCpXUYm763nIg2Yonoq6oimXcL62J/iOegjgjdWvrun+pwyysE8QyVl1rbXt7hDU5XR9
xqaxkS/P5e7Vs6OercIJYp6qQcgaMdATme/Jw7xJgsKkxg5nidaE0Cp8oBFQhDxiiKdjyGFmTE18
jjcyqPjr/Tm2r3g92rUNYx84+KqmDmhQE5UIC5IQO48Ekhxio6K8/DOsVRFn1URxEh98yzQWRlM5
egiZS9JMSI6kHadChkNblOI8/SDaFT7zc0nwDI4s/vhY7K1WQVxaKELWeiysGKhy5r+qb3GHgIwW
GrqUlOelfG8Bb+CFw2l8XkwA6U53wDQ/xBIb8Lyl8yt4gln6R31B8IkpgqItiyNTq/M2hpDGKIvB
PcLDbBYS+jdyuEYgTen6fhxMS/YWVfF7G3zV358XRx78wP5NRlwgLUwTbFtvWNTsnuqYs7ykhB22
qtDsy7hf+JjZ+YhWkv+oLD1EI7sUgRUIhO7xxjbX9Vou5mojBN4+U49iFi1PUoPNqf3jJcEKXZdr
fbnpfV0WwrYVnZ87xS/q5G7SYezqscRXhKh4gmJeemWyjT8k/HQjeiCKTteObsBSae22hiMh9WdN
lP8kNjJE20ou9LNJYwlUtQYIvjwdpNKkHfT5PYsI5xQZIcNAc/ENeawqcPxJitYSX1ZmmPMcZqBe
jA6TmOQhMP8hyqukGSQk3OaTX+kpMTZKW0Q+2GhCiYFtERYi6wkf3vFAG2sUuyrjKPxnmfLbuinS
viDQfXOJ8/3P9afmoYPPxJt3J2Aei/KJlWCC9IKyEViRy9+RmoohmjcXDJf9HxIqAaAT8BgmgkzM
EF3+j7JqjrSalXv+Yz/YLlFPy2CGPDC7Cax6HEl5yzB2jGrwrrQIjKYjJRwMr7zzyAHfw5QuLvMv
kq8EUv6OfMFLfVYLe9+Xupv2FRJ3t7w7DMCmnjCQP4tEHd3b99KXGlwyEWmWsyB14+QjSD1vxizm
Os6UuciZQ+bYauPg8I0nvzUmjK0ufQtZDACjFbbfIutNjYZqGsX+yWbyskOJPHLEeejuggz27lWk
qElNUqeeRchc8XXno35b2pOSFcb4GOWDTf+k7UD+c1HdpVamE5OJZqeXzBDvbULI1c8TxVUhN+e7
odKFJAbDXnie2D2ECyE82HgCH/jLa8I5HRoasmfLwgjylo1RXgnIe7zFJqttswQhEPmu46/KSadK
RjeVfJK/fbezQlYpi/2TLdOTITEMLRaLMXiat0RtjA42xsTgoQDzNA69en9mMq9OYhDed4YP1MDy
BH2DR+a4759mGWmRlQ9wL/5P2PFLTkaeWECDBfd20gyYExMNOTvqHG4cYdV71FYTWN5sQfkSB5to
kTIyYdsWfn3k3fD+A5oQD43lqg6ZfCzRsJYK39nMDusb4Tj2xztsJ64ZBMONgDKQ9D8aeAPcUOr8
EeXrsGXC0gkt9A4zvs19mWhCB7jjFysqVdm7feJcN5NN2+SM5H3IPah5jtxupe1EtM3eygNHiGdj
QsSVqASuv2hDRmR6ag1YztTgwgsSaOKMuMBO2JKgLI/A7M/LfT8S9vyJV5Quxh3fE8JUa6HjhoFB
X6zhQOGz5IU+Y5v/eCrhinZwPpc+gU3ymLH+djyZlEnPlI0+eTqaf/VsGhT34AnVGO0YnmTfjRpk
m/mRq2kXiqrAFRwxQxYkgm3XJrCTfSesj/FsFATPhbezItHqEyEcBIj7CiR76l8n6/UpxIaGcBQa
y48K9/YLT6SGpSeUYPUUPL3FWBP+WpaZvU+ik38p+e5Q7Jow2JOF7SCdAE2K/nMOaSGRtbVAZuMr
JTjWkvK4P0vde/SmjTyPr614jZ6j76hGc0x2Ye2+lGRtpDA2K7WgqmTe+ps738L0oqihzOgltOWZ
/TzHOtJbt0mrH5NQ0nWD8Vrgh9fFTT21HWPP+RDb4MxdLwWFwVHXZHl/GiOLO7+t3T4epCJsT8F1
xR+jXuiIPx0Md6ukVA7uNr0Sl10RLi/4Anp9wxgls3IHs7vTNNwvUZ5PV38zv4nyzDdg3aXXP1KD
S8UVZi71HeuSf8Z7K9pm+P9VrZ/gnXOu9B9yGdjPKUHkYJ2pV7u9VQWglfeaz+QdVbsvnTwseEsj
R/QDVOvX3Yj8LeLyd6kL5h60xd4ifwcXLdIXN3pkjQbtFJv7GE+1M8jEozLjDJ7O9HaI61BJWO5e
ct9mv0JCsSnDR46KXh5p7fyO9RZcwZhGYgnTaYOd9DycD1I4Dpm2mx54DjyaZPOpToUyOzdW/VeC
p/2CvxKq7rdZ9sZMbYVJXTP40wbQKgixHHAP0XoVDy1vs7G6kUsu78FsfJVbzNDWjaH6wwLgSx8N
+MCzUOaVv3QPSUIO3qpxq8lPiPiuiwUDLN49tme4cRgeJY09OVNdLq2VdKtUSiYOfzDz8Dk2ujgN
AIQc/4XPlRBQ2VPyKRqnV1ZIcEblsIXB1xxGOWGQYL4RZOZB8UTCHhNRXtkn8SBJGNcfwNhpLj8d
YwrkgRzD7/wlndi2L0mhQ34TSV1A3Omwefebi+wgpuqWp47FYi+xTn23Q9vqmicJVb6/Uk/KYqFS
q8KTh0uEsY+fTyaySBKDXDRQpJQ0AQwv2EWy8yF35Sl4XJRRJG/EMWltEYcZXpQp6or3TnsXNV7M
K9q3kCnR52IPcZYIk/1SvJhwZ7fhGW6DSYLDRKHwhjRoYch9sTL4Eke6yGj/ujIKFpu3fRFgdTj8
9yXrHLwzU7IVZaXxdhuzaArBqFMQ8UtcM843ofuaxbPvRN94Gxp28AURTIlocZExMCv/YqOqVGVr
FWRz/Ld5PfyKvmJEcO9Tb17OtSJzfVMXXdE/Y3TrhximRPSqdMjdjrZtA/zb6JdtJL/BTqNYHy5m
wzDSGqQAsrmdi0vOX/huErf/57xqoBh+iRD5mNmkLiQcoYiqr2dN00cxAiKKPWyM6IE8D9HmKNar
QiSFlRyPewSIONgcUiMbhwt0puWxwSnHqa00+2xd7FtTzMKitf7HeuX6TWMh+qFNgG235Ot/1ET9
UShtVOiEOxV/wIeIbuzrYQ+8h6DWgLzFpZ5hmrPxJiKDgxow0BBhu/T6nPNB6t83hYZp8zOm5MCu
nBkgNkh09GwUCGiOICLmjSaAapZj69BPlLX9TQUc/D3Lt+ydOGAQqv2t/+Vg+40AtM4IDyM1R2bz
pEiQ3+5rfkvbSeKFpWqF7kTT3+qUFHFMVbicSKFzaaer+OXnyEG1D7UiCylwItRbDL54mhcpE0uU
tK2+oIpye30HaJCIGknGM5igxTfUpmsDEhEoxLVokIQWLFOjR4LT0S7xNy77y9z63rcnCl6GEcwu
D/Ff/VBJxhbQ5L7AXZwTEQ2r9slqjsth/S7gH9lsCMz6OCCWuUAgV0D5UgKylwZj0k7Z0jRKXJnZ
XGuDFragRkdzU+HxDqDQr3u8ec4CD6fXxD9ArQWxVQQRZKYWVugx4f2Q7aeeOrnlJzO4UxPenqap
DfwLhGeHa9tUo8rteRLAA7Woz7tkJHMdNztzYcjC39NG85flTqsHOPy7nzc9awWJmfgu64FFT6/h
yieCTy+Mo58nHpDGE5BOqN/UFmngQfj3ppSV0Kpy1vYQg+5VxI5typVW25GRzdx+pPKOZ7mpXJHR
xj3zFMxtpidjq1yZISnSY8cHINkQMDQvxadGNTqcO0aKS8rPGS7zngM0ysLNWo4wJjUAhU2BK5iO
I/C/Sq+Ie1PBLRoh/tzK5YWoGTtlEA9K0hKruXzrR7tzyf6CqelpfhRuSsMwFfRK/ADYc8dV/3x4
sP9xVCepYkrO/K7N58Pe8f25JWmQvYtK3kbqbonpgLvJPboNPrrYfCiOkCbvkzJ8mmtLgIzqzigY
/BjqHvrpsaGjc/KWAOXOcbjUEeCt8yR+qOScBM3zLLVibgNbwp2NBQikN+SY2ShxCPTM8oOmQ19g
qafIazHC5N+c0UnyQeJOwIZccPNXFy3o/CBkOG+/AdnqYngMhNk6M31+FCaDEe6Pqi4oidAy8gzW
Pu6b8/xKk5aPOlul0h36AxK3apFTPkXXr73TVXbNtqtzGmqDKnIHGuBx4fFeyGysh0foxIdK3hYl
Pqa1QtLDraptcAcDFKHUfDRzTdtxK3kBFRJdKl2ja6gm53tD+ZlcpnCZT+uHZFDK4NiCd9Kb4eow
4pgK3HzHlu7Ycu+VAGt1+c47xrUjTMINoVWE/I1UyuCYs43qOil4Jvu3HOhiMko4Vzhn8l2qoW47
ND8nVXRvp7olM8MWJoboPKwu6CmGo7acDLs0L9OFBS2HF9gnsnxeb7+zy8VvfUO8WriGHL1jgAGm
XGPl7ZsQvPoY/I1ZOW2VQ4X7C3HLqsHT+DNojnVKqlomXBKuheC2vzovkq3nAwH2bKm3pLbYIx5a
Mbf9kVttN3zjPD5f5EtQ1DGQgs++EfRJ8BgX8uJqOkN3WOvSYSYHKCPR3PL3lqpiPqKvVcO0uOQ3
DaZGGSeomG9svM6NrbC1CAGHHgRYQwye2iXc4JnXaWBe7a5uRnJSNdklQlRJW7+1nn7KJfP6A0TV
XksvWi+i5mZOTOG4o1tgqueeq+ppIN+yHVn14GZgkbGEZcAbZkb73wc4Y1sHyGSd4Pi9YL4HRprW
81NqIpWZL24LplICHnwKvmsZm3A3NTaA/YgNOpo58dCkZ6/NBOP0KnxnH02aqQhNqyQwdAAwzFdL
tFTi9w2ijmLwnNn+2GnlkA309cUrjc1BqsEQZtjg6NjmAzxQPvNuYZKtlaixi2bF0vaz0UMjhCqa
kpIcqB5cF5iUTbLWlY+WcfYap4L0dCGyq7e4XhFW29shj+fFmUbETiOKYavciyX0dwES6T2QE7IS
MWD9kjyBWovTpzMKy78+p5eKNNZ7onzYS597JIq8f+O9Ack/7psVA7MPj9fLnq8iHeZ6NfwS0CIy
QWtclap13bx1OWcRnmoXrf9tShRAt/A+fhOMgCBmBATwviEgkxlLkBQcn2y+U/WuMwTucSoOPXLh
q/iL/HhWRG3luDpUIJ35d0PdoHQJ9khVCqE91MZSUAXC5egcNy8V83cBg+nfkFLmWzdeVED0kkxO
lKVBMO1r0A/cwLuDz57lr5CCQrdmJ4319m/L7JqD1aI1litBvCaLLalZ+115krQByT0NrFrcN9KV
pC1NB7yVtN1tEKQXs7jmE0OvVI3ZaeCjv8Ndd3DjOKUlmxkaavBlYCLwWDZe5N7HPmp69Fnrt0fQ
trVpVEmRkTLljFVCSjV4jv7EroxNN75/wtvimRbMZv9VvBVLWc7jBQPNJiXkph7c6OYNOXTfSDEK
yVnlz9qYLQp1gxqFpBnAwNxcMoQjpPwLoBiJzLN756Ij1kvVh3geJE4LyxYXLM/I76qRNmCA0NcG
64r9/f5fylqcMSp7pDt3AIE7l0XHsJSYF5cvkPBv0ZFRvHrtr5BpJUHPyEQ10+dOi4DACjY4hBbh
9wN/da4sh2K74uFk5XX4C38UnQobI+WytY5vByKwtyN1TnLzY3Jx4VptuQp7c7cFDx6uYBgQI0WI
B4cy9uLXqtG8PAtXgN3zQ4ZbOWk5+z0VdGPLae7UOLJo8Xeve7q0rwHsW4u2kcnFlRefoFtUsyxE
CvAloHR6B366Txd/b40IUXZxuPaQTvd6WvJxSN6z3PWG6KND/msRw7igvEo0qKNZalGVd7j8xfn4
fAaxEIkatGzPyNTPGt6UqAhBeq6LH2TOubTQH1BQDzecbzxKh+2+O+oNwOlOHbAjUsJHYE8oBs85
b6OxfSJ7GmrAsGHLUSAkNjAo7YZ9rFisiRZlh9l9W38CLFzrGd13jvzVmlGWkuM5U7ck4w0NSPFz
MqikSjT58nZpVPdMMMr1c20CIB3C/rgt2QzsC6U+oiwbO3PEyX8xEVntazkG8zjukSmviKJsA4Hz
IJ5s9d3jMz+8qWUHMe37IzsFux6Gjag+uZ0yflQhyTxtli8KiNa7n27wW4FmayD+wCSIMesw9LEP
JmtJ0GHxDfsymL6bGk8zWv4hZjnRJO0DMX5bZFTwGyhABVvhBIojBJ09Bb37Pspl6cLldwT8nTUp
OUN7L+R5ujEUk86Js7218ar+FAuIfTfOld5BUCJ2KWV3AL7xO2zjPtU1HegB08la0R1+s6lmciKG
yHIQFlaHmzJ0T9Asg3k//t2VH6OHnVTgWwWOGVRS1Za5FKni3ltDVnQscBNUcBwcOzFxLob5XrPE
BJCPd8jBfktjPWWNrW/v+QlXOdKcwvpL9yEI7d/3Ybq0H2rBOLbu6Fb6yEY7pid+aj2uw90pyysb
B99jITf7EvIQxwQZirZRqpMM6JyamFZ8p93qeBq2GsLBL15ey6TbcOFe33fw0MCaOsZKY2TE2ozT
AFq3iJhbQD9x9rkHvvGqV+Cm7kjkjJUm4k2qxihOCci9R8AgwVg7KJ6pCnC4Za8sX0oBQGg5Kszs
z70XG+Vvbwvhc0OWoFbiyt2ViHq2EoipVlqauI3e3g3Sl7a05jHt4jYvVFYfW4t7hdBDRPnN5ylg
6DmTRTqY+E/7b9zk4IFag31QucvCAnwt0McF0ROTpQvWf3mA9XeSUdTJmz9gBXdYe2koAVGE81yv
PFqhfvv087/AdqvLpD8rcsQFIqu6czNQBjzGznZ6y2QBO4PyncfghbLQt0lnGvCJ+7KQOvmfsswM
BvbNWtUZWxHaekU8yevrU6QuDYOYXbXphGkoPwUks13wbqAx/RThdfq1j5UcPcN78++ue8t1majr
CTYzVfcxcuBf1kkTdALAbKH6pmPObgk7BPT4A+jWCD1NPFdKDwR3MIYgRM8ekqNf7Ab+M5V26BVV
5IkvUCzk1CShdWMvFAzmr2VqWg/1hDOuPdxC+SCXdiJRAiwT7OqXBW8ZVwnlxg/F8914mhA4CgBt
ujGlCXouBOPQcsBvw9yfhxteoC0l7AJ/1QBa/bqCuClMEc/QJyBkF7PMPY+Y6JDfwiHaAyAR+flG
uM65X5+OI9WmK1LH9EJS9TuK6DQgLs4/ey2SSww49vdzCN1CvSIEa3FnUatzWWlnUsE97t3Z3jKl
bpcy0XruzCUwCB/uW26lA00Hz6Q+GnWc8T6FGrVTsH9v40sJxe4FGg/LhRX0fExwRaarZo23bm1b
A0cxwJGePcSbUdFCCacMX//vzGv4jO9ANbfoyDTz3BBSjsSmHBQpI/vDogpBjQsOjzOxCumGTOiK
aUhnJ6Me59LRWXT+1Oh5qwUj5MjBlKDIdT43s3Kyms9Q27oFDYs6CrDggat5OjVH9t4EbMe2pgA6
XFa/n4iwgznLMYII639wfH6CDSrkncgXE5MH/P2E5T0OcX8jWRnyx0xdsQsl2e7p+qdy2cKF0NlH
XqD/Jt/19LU5M4YM/xkAWPWclQtFL00YFSdc150jQhfvm0XlTrl0sHThVZcVQa5VuAMk240ZQyXS
1mOSBfNrSk8rEo8yNfxM//co9pqDKBtRjz7R/UtuIFZFpW9R/UiAD0Tp3HYfVfB+IaNGJpVi3bDt
Xy18eFY2A6qXBRf9rb09L0zBLOizCa+Z7+4t0XtF6D+k3rpCzBHawLEcv/kUALfjiFHTA71Wkx2x
CYwLzJZNBLAtEnuMEnoKSpOrzD11NqniS3eBkKlct1aAask0VyF6YR1+GPZxnN76JhQeWHTJVLG3
06QwEjWseTdZu4hdZahAGwRYOALOdqhPgM/sHYC3qpTSaqSz3AcxItQkMfYCXFANryPqBckbeDmw
izTC0fpwvTO/I33fDAaRSGrYdEH343JKJmO80H8rLJmJTWB3B40tRdPd2PQSMzDYHLQSiJQQscze
x/vMJzM6c+sfSuyaUngyzgasaUUcSdAEdEuoZIaI8cwYq1+WARZm2DszLQwqnH22rVnU4ijS7J7I
DdAgfG3n0MgUIE4/RtwVghbOEX2AFWTXtVBb67W5p5dOM1BW7pTZis8BHoOzkqzpjsG2OoSwgO/0
uwo+xKDH9LJWQlF7r16A+or6bWCAsJn0MfX/ImPq1Uyk+iaiLnfo64oUPKC1DAUnx1cbTC11Npg4
yrNZLsvdAss8Bhytej2QLcucyxhKj4AZcrZ9WGjcQmMvfx6hRKsqpcPLJI1EU3gq7/k4gaeDu4/h
yuaixsriCcd/tY8Bp/S0hm1B7gZDfIHG7Fs4Bkqm7WRrTmoHCwLQ+4Q8rB5NN/1H2WwJOdlQgp9N
6VTcsZhkz0bqZYRe6AgcGke8cuB0lV9ZFq5NjqwFhVn/6U69fLrMQD5K0xomosqGZMt1SyXxuJfS
ldsDFIMf6ZGBgHnoP/Yelr9DL8BHeGh6ncjQs/ggxlqZOr7PcQ4NE4NAh0Rx+Tu7rDtFHtjSNeCI
/cFYbuYSRrQKs74Vz57XkrYj2kh7NBGZDT610B+bu/0h8Jya840ag8ar8DK7CE/TYNRr5B0jFAs9
+nrVcYXxSmSBAY5OSoAUU896TwoJKSFvkNIpbF7aA5ax0xgTI9GqZ6CMUxe/7Co1Kfev5UNpVBqt
fK1faD+TZ4dDYByRE66M1lI8vdLij8kGfJQxOS+Omb/R51ibdVNkWBHD30/e63aah45OrFAzDvSu
56iPzxIlFoT+CF20GCzVkIZU4iiniNK3MZM3dKH/uU6UMiGtxc5JnGcpsWlp9bezDs8AORKoInTa
ckMtQHJjgBOCByJhO2UcYLy4lWO6tjnd3RTXvWgDUGnJBhCBMWG+a/F8qrxcKcLu/M8B0xKacxCo
hOVkW+aBRCGPXp5GpSO7gRyyyGL0zbCTnUNA2leoOyFJ1Z/Ty6u4MYhz2yMXA4iims3SO8z3P6wX
KVwGNb+mnev9ot17w7zRNFy9iJEJRj7ZVbU1O1eAfbbyv9MBTG89NENhRem2/2BaPR72ye9xO2D9
K84ksAqVSRXnUm/JzKFF74LyHQN1ecMdgwdq5Z5nLS5n8LEp4coD/ilaVSTe98AzzWy181cgxqci
K6RxQ5kgjriv675yZy6RUtCG0CthAFzaFIzM3Sk7mQsXSuPolP6zImPFXiTNEx6gpKgJvKbQac3K
eE6RhmHUsMNS3Wp4knBtzeYtsoezYaUSSvPsRxN+g/iGRxSynYZzwLa7DLr6ATaJPHi408Km6+ez
uozYBgbZJV2U9Tg4xcIQtZWB+kArLd5klIXtViGFW7Ki4/rJ7yVLkw+O5E0W8Ll0f5w7ygF1C6Gn
XCQnvksH6Y3gXAev4JPuLovNzxSrsUMh+br9qhIVgLKXCqiDvvDHAALTNfE5LuhV4UGQ9Nx1QpDW
3fyBdc+4SRCGYFUAfbyx7a+f7W73dyRlHEmRijaM43eEtBbbojxzm8697q+1Je8BidRzdIqCxHf0
trja7yjPK7J7trM/kmZjybSb2Ohpcej96EHr0/iKy8vhUdQcRzuU04z3xW9nMisFKlkufljIEAgI
J6QlXjipFyxe/6cAt5cSIg9/xLe8yIY7Hf5hpm0qIGgmiwUF16Owp1ZP+IoxjPcdU7lNK/ELqUz2
LVveXULhnCFTCKNZNZbTA2ber+nYFt8Kt4DqxFEIv5qKIngGFQ4TI+gd3sF2Hp0YfmAoOuBfYUAv
WYeuZRRGzz982L5nNjF40yLB43uIRFFS9bfg2DK1tQpQfINku4Na6oRpY1WsdChqPPYl/CsdRIy9
wnS9aOCiGEHGo4RXNjkZLVf1I1Fk2Zrvfe+VtCB5wNHqnizhvwYBsz5io1QmLBE8LG5kUjxs5j4c
SNscURoitOWpQ6rrBkH1jHz0H81h8gjaQ+lUozp3MR7Dme747IyxM51JZSEP1Y3pb76zPQvUPSrR
Rv33ZIAJ5Me9OcqG7DyFMed2xvpMjAJ5JRWrUjORsDllR947alsGf4jx/JsoFIPoN3k5PPvc4o8H
k/+UhQZImYSudN5gYRjXnp5GeiVE4x0YcDi+u2T3Ks4EC7J6kdoTMYdGRrlX9+fOt7MQQgduCpy8
GeiW94eIUrhOJihcMuq/A0ueT42NxMspWi0k4oVudkIYy8CVfz7cWtgLsAahaY/ElTpXrhKwddDo
s1ioCVgN/wufKgmVKYaNit6n+WtQbyoFdRgfrDlFn8fWInG/xda+G5HD1zsRDbVJhqHWpQiMtLyc
yYp+G1r4TjRueCVgwUzU9vhLWIgp4yP7PWETHZx/sbxmWPyruOalzFRR58BPoO684zgkajMerVfJ
AZBxc8EeKo9IUqPmLkdZSPTUPWGIk50STze2+KmEDI6LME9gtpHpJfpEs4r46udkY+0S+CCgGIvz
x380ntnGA6ykgBqUR84Nn4U6Og5FOFWquxY4l+3AkTOCjtcjkGxkGTs/b4O7Epen9CX7j5PO6y5t
PxgE3KrBykHUH78maT4nk3IBk9iyR4CdVdbTh5t3mgfHea2YIyfPIDcSeuH1aVX7n+iXQSUGBxCX
Vb6r0W0s2LUjjeDNUXYsZwgYhzMbJT4ffZpm22k91cLASYvu0sAALwc2ArYK5xxR323V/YEiuIL7
rvGU62Pflyj1xQJrSgXuWPrgr7uh7kHZw94i2oNZ78mqX0eXJzzDsxWtMdowg4Y198Ok/m6qH3EA
1EIhI4s/lylGwNzVjRIflf6yf5aXPEUwP/ITvnYXwOk497LNQJ8J94MbjYS/mLrCprbbN/+hKWWW
OL2grOrH9Qw5bfPhXNa0dqS58ZNILrnxhwy21tZn7U7A4/W1OzDw/8L9HdCkQXfBSav6RWUMd9Wx
cWZulI0g/1z5wA7y7D8mnGk9ePacYEQLfr+wCAfCiNZsaZIL9ieC11fI3Mr6G+zF2xcx/e+a30PL
95+ovfnp1LMu6wfcFbKOnJH5dv6XiA2zFMQ14IEHVbaAwVTezRycXl94xq4zuA9aPVimF6yU+3mp
3I6BQ+B00evOENYnG1cscwbQ7NzkPar8IBiHIbv/mu+2kskmgxVZpmuEOgTC4F+EUId1v7mR8YO+
4GsdwaOht5xxRiMugjXLJesQjJzNUxOoRB9bCYDahVzwbPq451EBeI5XnagMJcBTV9BVrHiZAgA6
fbZfqvFUdcwRzqyAlSp5YSyspjO1/CCl05QYEo3llD7RDHibCOq1iNGSZRAc0tpG8uSbXs+CvBtU
Qm30VEC/fToIWTSP7QFhI4g9JqvCfI4/F9OvQLb6oOrh7KQ9cXIIxk4CiGZ5rag4rC0se0yxDxac
zwyE50HTetmVNv4XOJJ7DP4GxjjeQ6L/FXhYnrbz3xIc/nLKfjUxvWkTj25aWYkan6CLXAkU7cwf
Sxo22MVLqnXd9o7mhcbH2NIjeicY6fedbrmmBREn0kcF4SPMmbedo4nuKiw4Qa5E2qPlCAxDCRco
SkqhbewcQSflV3hqIIQYN9R9gQJKezYEKGCKR0otQxYZYoUDyhS8mSaoFv8sI4lZrygvePkIpTgX
2dCJFLkvawZxXbZHfiz6sea3YiPJA994bH5yD4c1OqFLRBwp9OnBfwwwZvpwi56eaQrx1LxWXqqT
Ve5nfui+knlbajtWouEN3/cLT2oDo0vb9wDUwM498VNhfvLDdbVLIAwakpO7LSu1/9U7eH2rw2/K
r3R9YsuOy3wPTiG0UfwqrL1OpLIEy128r6bYg8N2oiySBcs9xIZBg6a4rld4Y+0njT9HbHbi6Hxn
Nz78yo6cRacTUXGBtTdVnM7IbY+dptB/m2d6Qgkw70wZgLIvZTLTbY08jit06KBow6RZiEvcW7JJ
JCq72PTagL7uz+4wep0L2qIyF94hho0wTXP6VdZc9NyvmlmyckQDo6eGIUtxmQIzDhziyZd3inUZ
Tg9G8ycqfrIachnbKjEtTG9eKPEuO+lm2YuRnL545LuGcDpsIjXMBHQqlnoKVqOiurxqCTKYI8hl
NR+yb5UQGyKb/qY73q59TU0VXY4A4rzLAwOhmECTov/Ny7r5FNiMIPfDg4dNBzDj14ilBLwRymDn
9nVz7pL8kq0+LEemx1ImCGRveznG1QqgnCt7gWrXUNls/Roh1D01I9o1uffANnpb2Ds2c2ko7dxI
1cyqcNvNquDENCb9EqRLU+3Gv1dc7U9Gc00A5IIuf86Iv6baSmMAa00BHj28tcbqw2j1b8kt9bOV
xL5NT64liycwkvGDzWS4/ZkaV9kLI2UQ98m6a81VzF/ELBs4FCbmI5AV0TE0/ALigletJiSgOjZi
LmGKbS4168HKTNHbgXxIP+RNi/VK4YlkIfFq4/Jf9rJZmz/RW583Fv943PbazlbKtMLYbsd79D8D
FN1/TXG447civCa6Qklq3SSgLOj/vZnS2zcNJa4XXsuHsU78pAm9IUuMciDVY9RmTHi1MTo5agZ+
Yy+EQdD4aCv5reQjK2UwO3dLmlh+W9EH0yNELSqRS3eJFS+1945Bs13TTR2sNJQInVmr2cAeF73o
GfZZIe1XJj7eiKi97EwtWlnCSla94aAE3ZlttjVfejPfQlH8PU6T31Q8gB26AsfNHcPTvM/JhVN2
koPVD/MQ+awMCB6qdN6/eXrQgmayIpycAsNHOuDAyJmTU/E8YpYDHSwb4dahPg9MevtuRhdiEf3O
rz/tVlupES+M9YkJG9qUvGPz6t3NN2JHVIHs6MlszMZrl2nlPTjwacbu6DrX5klVsT/FFbxD1Ozv
5vrWBi8g8pgd94HTbhQrdb+2MIg7LWC8wIujq4OriOTja46c22u5fjCgEmqtRI2eqlIyW2mq/MaE
12ftXJX5/ePkfpth1q2Jln4cdrAC0YQ8ggL5at21QrW5+kp+xf6fxDqa74IX1U4i0WQXwubv/bDb
b5pOKz24Dp5bn3tVDGAx41vsMMiGOB0JDcZW5KNdNUA3q2BwXq70heWsydQKnjz4/qk8N52Ehsfq
y7elkfBV083kx0e7KnY/e0gyOVIDoGiZFRoDtOOTypSlCQrrrCZiFGN9bpq1OZBt9ryYZaN0lftx
u3NJxjUavJreJh/qb61Z+Jh2fIAp/NyzR24IpNRbhQC9BM5D/at7mgHUy3Wk7DxVm8BN24Kdnshv
ujaie3QDsIrFnVOPuX3xB6a7GH6FQp3mXMxrgGs3glUFEQwGG26oN5TfcvGE/3BJz5dES0uxmMle
/fRWiwjQaLHaG/+c4XKRZYOke7MOC7cgYJaDSjPjodUicYeLlx7S//BZo+l+Nr/AeU2x6K3WnTOp
9xc5Q3SX+XNrW69AEg05mlDTERoFaAm7/fzJZjzhw6i5SCEqwO5fj/kyyBa4GX7orqpXoAA/z4qv
o6VqgUbmAv/LIiXoE/u8mZydnIbbSWoaCLK8Yfy8/woPmyXCcVEATv+MgVjGGnSG3nJNRSV0x7pV
Arscl5K58KnlXw5+6jSal1f8aWA7UWboF34EUzgAmCxbIhbcSwUFB0xFVwPdFz3kGrKoz2vKEl98
CAAo6cYfnLmkRaede9TpFMWZ/zwAugegu+o7+PDsqA23IDXc1TFLeb7DXmGWctjH6ksV06PWCJsY
Z8I7o2h7udK+mCDKYXGxxOvkyvGcvkV+JJKxUI+n8mkwQjEYwLhRe+NG4aKu0qsv3gIiyfgM2Feb
lOL9ZAvJcX0Xhmnw4MLM7fAWy4hN3Eg1kpuITJeb0mwhFKjRMs7nMLOG27IznoSJENgkOQf5OqPb
4/TZsmV07WWkeNmMM9Xr5PglFSedCMEII5P6fjosv+Zm1vpcWgc3185DuzbHqo8ss40p2hon1Ixk
V6pFF+xzSgtXcuKe3i3eA9B3Mqea8qQ8rSZ7PSzefpN7OH2NVcRiW39eWsBZdjudeoeNytAWq7Tr
lTpp5NKB/Tvog+qhE1GIYr8kqJM91DazXeF4/0+XIfS7S8FLLfqYgJs6P/6Fvi8AW56pucs6klcs
CaJkNZU9EG3EJvtKU0xTctNP9jZSxJlIle5UsMuigczbjU9ZWKeVTuPnaJRYDJz0E3APYxoBb6ha
1+Rk2/lhBLqezCOEhMRNSSzvE4yLX6shLscT+w4pszhwQIKWOEQuCfnXWPYZG97fdJ/29vlpBBQI
Cw3ZpAYjk4DAyVtr9aG8GJZlvx8ZDJr70OIQsnhSzl8tRwXZ5dLlNzMpkHMClmaAhWRsC4k0wTM8
6qjwQHgLsJUid/PZLA5xMp76YKoDLNPiHoSDW/bbnMimeXEKcHbmd4HSFTrQWa0LXq3sQ+6kmEIc
zvKhWHf+fjL3SAD9PLDxAPVBxBVpDciX2TxTbS/EiE+uKbLPHif1kmzFIbZa2ciMYr8ZNuGpcsSC
rn1bdnGoShIx2Zp01Kp5TdR7UF8Lb6sZ+fKXshCnhSkKky9P0t9Xerfgk9pFn/DkEhNb3Wg37QEu
cJtsLyB5O793SLhMfG8C3fX5X7usnizidgxafC83NhuWWrf61h5p8FKnXR3KZcsCriXy+ZDFr39x
boi/S5hbA1YHydGjcUmVJ3Cd4Fsj4g4iEhXcoU2LDaph2OK0XW9I4WDvRBOXoiIKV1Ywjc3TSeg0
hsldseU/ERJjHK160V+bvU/vepE8ysAg06/sP2g5A+7d0t28hnxJ3uEiqyqPSqEiDhSF5S/hMWgD
eUz3uf3rfC0EOfhA+f9HPhorTQKXCtRppWyDCYBJqBvEJrgZOCLZKUy6GRsjPfPdwcPcNb9CQ7Yl
J8MFzuejDg2IeOxJ7bSosZFrSbKAYZa9B/bvFEEDujKPAVhvAhILDgggNQigpllv8kerQzdVeaVV
7miYlBMK06xofR03P6imSNfMdWDcgbDKAkiE3SMMJwhyoNYQu4844ZE5+rbjMO1Tx/uOr4VckT/l
2LJZ5FnaoSqdPfJNtbSAjdYjOfz9d5Hn0crwuqY51ECKANf2uBo4XN4ZidaIn1EYDGkTmlzla8D7
o2tMHcIR7a1XBmn6pX9yb2tBjjxCtkJuhDC7f4def16W4Jwr2fLd2YnqgT8PnWMtp5Y9nlWz9aCp
aJ5PX14wsxiteujQLhK7b/59JIwjHmtZed33MC7RgRc1VOOvKIwFaNUmZCwCjZmcM4QzkJUJcgbA
HkOasqz7+hCn2j/c8oYqHqTHq9eD+VMFxbYjJ9QIsYoWNtS3Xoat5YIoZEq0liuvV+/wAUlGuMRY
zz8DSz2FBsFhZmbRxuiKZ6irNw14IdSjGp8tMKxUl7R99aMfmqgtJwFES5eQVYOGltbOHLGEqjre
ukCdeUUuEQ/WJGqb7Z/00S6WvY5aYZ+LccFPCtElNtngbkfwikxE0zOPSV81KtmgiC3qNF9bf76/
6GlUcWKuGYf1YUgC9RYphNrDwrRPHUwYWYKtjjrqzQnA+2KT+TBg2lJ3LiZt48FFWyC7C45J0oLV
uux2En2q9XKX/pIJ5oLAn+LteHQaKE+hlp79mEq2sNp8tScSYJr9jQ0ftVpMOnLiRY9Ik6BQAwxo
KS8wQJGRYve7QrF5VttfBmkr8bOuRwg6wwAH8X1v86bpN41eYUy5XqEhSvVCIqxM5whS0AkVErU/
J861RH8LR2gc1m/6rP7+6Or2Prew9WSBdISTMGzZ3f4O7VEw3CQb7bwxh11WIeeOyIw0O9UTo9nE
Y3ztSkelbWTVzRYPfqIbg6UXB5uAAjX1681W15uukhmn2M67NxZskIhJrrVrvmkraZYAdXrUcRZ9
N0S1wmeUpUn3BS7YvJx0ernmMLjUXwYuZgKVrZ7LBFC2YbzHS5MFFq50VzcW/TLOVFaLeBSiAfaM
7yvXiKsv13lZoDtA/ELF6l1DX9J9Kab1BUkNIjsG0PFmGQlPEqDsIgrF3irRGqFBIk7KAvu6uGl6
jR3nXMRIn9Kps1APkXeobhnCFzKLZc2obcNWvfNtngCML3OXkXBYJDuajKJECueC9GjrdgSwcZpy
Mh2FYpshpF6/o4IDqgphR1JxX351tmqcgztHi6YJNFXiRTjfi9UKqbFRnESADQE+8dKSVJXby+fq
Zj4iAU4ZSpuTiuGCNyUKv9Sc1dtryoV4h82VmgJRJdEILJ7z8+u+niXLWuqrpf9BQ3REKe/NbDQN
crrrK2NLn8JL4lJq9+cpNuIqAhmWhMl2uAXtchy6fS3pYadDMBSng0sl7m/z5jKPXTnKEzG8d/b5
Ka/HKVkYhomj6/w7FZVluzRxxpbxaqRnN3JdJTanUdDcLRBjhu+LgfKToJUnW7Wkw8Ocwk4sSWYA
HavvYGwa21JEeQBCg/Kv18b/WhQ/0+lVM/BR8TbxolQjWpbIdQn3EwygKmEGbLweBMYur7npawmE
LGzUylTRyfhALkvjDwz8qisSQTup4QjQXP4kgWxbaoHc8o4f3qytHmM4fiw2TpL52o4IVrWqtYJM
bAskbn0RlNKN3IlZprHWmAu7SfvV4GlQImeWGBvc061vZYvRUDXrmKbKgq6Tm3nq2yJIBU8Tp18b
i/HYby+7+CUUsoM+MTtznbaefYV1oMOJ4DPYEXGJZn5INOEn7d/igrzaeZIROZWG+schUw9GdyTy
g8rCOdldeonDMPLxH7U91IDoIpzQZQF3JZVgWTNsAan0gBoHUgxnJwH2onEBf53WR49tD6nKakMp
oPBAEVRYLoj3OoeRDi0qYlH7mAgkhmPQyQS6G6qW1QtvrXOMbPqNg1bSWRwoAY1M/9gQHbQkzmWO
DWuWbZ3Du1gVhiKNTbPjbF0o50F3hcCFiArSLxHnsHnMyqzP1KyKjB7zEAqrNpqvtBMMyLSxAO5T
gpYmAHlnb8SSAKCdGkjKViCrBq9LUnaBgP53/zdub1zlZf2RUmClK8mU+osCVGUYcQopsDDn7uGc
1RSw1Zqzjcsg0xqe1HOwXiGq+SmFxJkLoqiJwIoeG7zFwEzw0bn1HYdPCIUtkoEytTvb1r8dwhNR
v4rNlII1Q/4jIcXNjsn/xKgBZWlyJ/t7BZU5duQgvv7vLyyB6Rf07FMoJtQd2Mo8POKznJuO3iqf
iUE6oOOmrI7xUjuTyD5GhwTIdUOmUGxbPvQBjhz9HD40ZzBU6AhfBkSR9m06lH8ab51eaFCCOTdx
n8wEy3px13T10AsgXqptWrJ2Bsgf6UZ8BvHvpy0dxMFGnlCFm5AE5lHm0V6kcB8v4SQDEzgW+f2j
5Dj8tQy7FsZUlqllevol+brWJYhiiTHznsiOLIiOoGfE5U59mVkdtUJbVfbt/fj0QPHQuDTngunR
xDPvz0cJvBF+KW38hnToFAUwv17xkUSNvr+Tm9411gWVoynwGYmbjX21jmnR7jJqWaO6e+2NwA9G
0rDVk3OPnpNc+OM6iYySzd7TytkL4Se8D6XAmv/06+AgPGfRsLMn6CYtTiPqHc33oO/Q08s7OY81
YH0U/BHpAX2F5uYNiLnLkXaEjUoiTQ6hFj2OSVWm5wcZtPATAkpOJvea0EsrHy04OP35b0SdiVyx
tOJ11EXaMqwgTdPgx1rPGYdN2WF3tJnpL2cvi6XyPPhDJPdiB44tW7vSuA1ZBJxbSpMVmvPru6Oo
J2uWbKUp5V3IKwHl80B9e1CLiU6icLCa/dM/NjNct7+qseM6IiLzQdpWiRSxbAYVU+khKi/QQN+r
jBlAznjSZbwGykR+FVwRJEuhItWeEi3uL2wrLz/rnSS2uduBEzu04jCrHfxwvN3LlRF+BX5JCPQG
3YDGtLVoF7I5W9jtqDssrpz8q5oJhHfkx1i6XhVlGXc1gfykqrOMK55wD1bOANJ98Dpizdceia4p
lO5CSOpSQ1A9j4mO9mUSbt/2t1MXNx/Pdmldblgbvw288qDanMeoP8zg4fvGu7I5sWZcGdHsuWYm
3wYT1sL913S+Z3eCF2EvfRjm66gzw2Y1wKJqmB0gyQupHyJAknzMnyYcLe8780uFFlyRqhjbRYQz
Nnw1b0Y9p04ll1nhQGoNdO29ORivhtx+E/HMkzBni67nriGTN/adf/Evdyh/sqWRtdPk2QRJVTPx
Gf21swX/3TbbhoR7zaEm64DrXno+K8EEc32y2FCtoG2XSn2nvnUtfo12BEpzzEAsSBoBO8EmIryV
5QRDZii64DETUmdW1V18jkPFI1jBdqUWBX2qXT/xIeva+0nL0X4eaVll6QlD5PKVg94FlNeQ922s
X4KQmuMO5admNSRitWyc80535roHLqdcdZoUeIW6p+EKlqrw5ZqbvTbbUayfJ4L9IksPHwr+twdT
aU4zf+7E15MyraL5GToVIawwVlihwavPZo/htyk1o0Y8wuYFKMi2NvPOeAMtNjSNLKxg37k2pUr4
DfvUGlLuqzUnHkQ5myrmUeKS/1imnZxqRTPhQz1xZIFsC2dY5nNM0IseO8xWdqqT2c8PqZ0/EU8f
/gQwZxA2oKVe/SacRx3HSqCHKzPhD0MZw8XqmDO3vQFbT2XWah1tDcfCv7Q0YRtyH8hc2ok3EX11
3VmTgNDCCH83XnDgTByqtVrbSvBafksn3yfeIxO6L1URKMeen1w5teujlxiwm7rHzwYAHoow4JW1
J9SGkXe6QXAL4H1RUEA+/tt1fEr9HvJeIZZ/DtoiBAylk5NnOxKyDCQtMUh3FQRbaUBI9Z7Hq70Z
dn481i9y2K3PVk0KoUtZZVN6RaRNSm7NHOH33wOoJU+vx2jJOsZR5mwAsrFNW2+UgpZzBpQbF7sD
NOYNUOmZf/0bEaw6VWi+bTScj2p6mgpHuF3c6aEAtekKmPM0nsySIGx0KZN7cvJeyZ8atzuDkqTt
EKXiGQiXA2wAJ2/qL2jX1yVnpPI+OIuLY2RowOTZIFv9W7Eh7jOJ+WijwsYX/3Gig517bFBQYZUj
n6PJs9yf2wsXYxrzX0NXZXtvPDBk5/VbpASBApw8T7mJclvjZEfqwzuHtR/NvM/sFfaBtQNe37p4
IgjzX17vojzq+Y2qtiRoKpev23ZiGq4Jl10FIKXdFXrktztsnJ0rRf1HlX8hC1Q7ODa+FUtiBzg0
sE4c/SizjeVsYKI8MIUMiPUNhHmgx80dltflRzctBO13AL0ORPhD/QO5/g2wmS8c/3nmvo5cDcZo
I4PLI1Gw7a/tL2SYuy58RifGgBrta9zawApJW7T8jVgl7lCQwtHeV8kUKP1G+JRkB5Q/UalutXeC
0BEzhNeVfkFM485MFUhja56EcFA3eFJJah0/cCvBQoHIDjtELVMUJWjfcJ9EXTCC53aZQlN2wzU+
kh53c+TFY/XztOG3o3ONke/G7Aw2YBu8rY2nzPQdAK4PXjLVq/pxprVjJzCIH9pfFGBoeDYEonTT
d8w2QLKXYqtewCRZg0R2xriSqofqwq780GW6m/pKKWvL3AsoGZ6dXkC2SaEN2sfGlAhhhbtjsgoG
/lNVXkAc6Oq3vK3eV+42/ti7IaJZvzUemVZdcy8DYRYPTPGeL4/9x4mM+TpdkUSVjBygqX42ROf1
NB1JfoW/gaPuhz1rAWmWLYY3LdatseogZ/Lv7TOLf1CEcTgOxpWIhemPGVSHbYzw81S2buBEN3Pg
IqHltbX8LJEUnDcVoarYC/lisv+z5j1bY832hf1O4MoaYE6UsoEuaovOi5LskbtIknW43JwIeH1x
5Y8StMP/Fq8IoIYzBgYgWKUtQusuuANcK3sZYTZJnJ16fN+eU6iWgUAeHSFoAWAEr43YC8Y6zszN
bKjIZTuZjsn8NMYsqPA0tInxkkPhixRIz1x3CnS8x4O/ZLz9hanQedAM0yNAnrkNPaSfHEcMcB6f
1aNHkHfipTMVryt7hAQ+wFZ8eDiaiRTQgBXVfUKcN9c5KOgTb25ohZ2SbKJ85ZeSKZqDkVqT3c7x
6oKu3vnR7BC0aC6ziGTAwcXXyrTRm2bMhfWwgbOgwMy1qIQ3H/c+Iwl5Mv6zml9eAL7opDPZUtvJ
4/SSnlB7LowO/2igOgMIcNnFINmPCw84j2GPcGOuB4XbRH/bflZhNVdygZ1gYKQ022/2kvZpqgO1
A2xx+3spmzN1X+Fcn7U95WvZOPz7ywDflVqOW02W96Oavi8k5W8VAYLNYAbnw+k+SBGiZJFC2X/l
1doXe4dBs63n0rrriwOIV23ePaDkwX5+gyOSkbMITCJw3JoFEn39sA7gHbq2uvp3pbay6t6EFc2P
FkrlifCHJOC4UGB4FpMu0HQAtIgbodyxnQAqS5l9sV40eIGeOEAn1jjvb6srRVi+sLCv4Kw78i+o
IAReMhST3tupsQh+8qH/Fb+3g6ehRKpwRvf9vx7ft4HXWBnf610Anz9cKe9fTbcoro97oJ3owtIY
UOEaSPT/qJ1fwAWm6b5b3km+Wh7OqyqDnBkFlqlI3VKy4M2sm80AKHMsKFTubNFGvRTKw9XNw23y
32pCzxGra7jk21Wc6jnJkBpzgKi9dAh8yB6odGr9gWRnHNyqoSi9Gfa4A/R+fwIShqFzYMHZcMgC
1Kvwo2tvo8lEsY2GmdL/AXRr+kH5UBBNqMdY4ceYkxiB3MVKWAMtNjGrm4V0EjUphmV5Bw17RlTJ
t8XptevbQbgdpjKCkqFR5mAueQafbO/eyAYCajRHhj+fNAzU9XBqVFnp9NmpVUEx2XqKtqkQG4T6
DKvVS9U9PJaS7M7Eq6c78anddzI9HVecYBm1DxdF54MvSX7gheFcDmZKQ2yHwExGRH4AdRTKEi+z
wbV81Pi2sK/o65PJWrOlQQGik4IlHFDqAidu4ODNjDr9um/xfBMqNg0b+yFyqiJMjrdGpx5zIcvW
Ov7mpxChKicAGiwxX+J237ddDXAPTSq3cw9QTU79qZ6kdp1Os+6NIkQlvH3FEpk3N0Dv9dcCmdoL
fPx8yyJb+tT1d5HrAJgXJxTESZ4qt7giUgOAjbNKc2mDib3vfi5H6/HZI53zSH9VT1gSYDoTR1Nu
tCU8qGOLLdJw+4hUcnFgpfd2rhIKPSYId9/4spIRwcmNixEFM/qGwOrq4qaWCj9hdFRCMh4WvugA
cFwSfkGpqdavgJzVYxHfciSNYQzZSG51pNJfscqIPpBMbgsV7hDsqPUo5K5je9LEqhHih4SDecsK
xBGx1kVwp11Yu8nsn9dJdA9YMYEzzaD1fKnbdmsNP3Tlm+BBfYxkCO3XkBxMOj3Ge8rS0T1zJ4Dv
xTOyx5/bx8ftc3A7pa9fo3ODOvYXL05tN1Rrnic8pl46iElA5QGaJTqVlKh5TfI5cOtcXg5lmyjm
Vu7vdbpi3YBPcCKD39fSKLkFpa+elq7uIDekEtzPcJV73nCi/AJ9doA9Hgll8EOdPgIBuSRzZk+G
yN6B3E9dFLzTSjiQGqGmZ/1ZpRZd/YZRbxGy6Sr+GKzKE8YbJszxfPXsu3oarKY9ewziNwCtvPiC
NMxh/okniu/Dl8mgtebwd06RWwsjBTGmEdG4S5MnYlgzFloY8WNxughAftCD9dwQpc8AJx4HPuaA
pjPNcpw6qneFnc5UGSS4oivNFAL63k4fOQZgmvbuewdTHo4hNRZaNxRql0aSw7yUSWDsd6WmmAur
aA+pRxvc0dBzlOv/+JKsEaUgQpXxg7tE0O6mU6u21vfX4LjHgq/nZPypk6aIy9IHNsWLUyHHtUHw
hGpdKpVA7whLLK3HfrxkqavzG9vyeuhSaRCzXrlfowdU0yY9cEcF/Jb1PQl0EHbw8QnGZvmtGJTz
Rclcf4AAsBmjQ5qvxT0D2PYe/SAydMIkwcB47KRfO53HBMR/56rf+n5AvkCA5r2Vh4IZ+5ci214f
4nKhp82bwePVHS8yelNvLFwOgqUqf4v/XZFr63OhZua2JIn3EdHX1IN9aRwRCKxGR6n5GEfDTO6/
V9wg/ea6hVkkLlC+Gj4HWyd8nr6zS4PJioOCGOdFAL8WHd1QSSLtVMBsuYyzxQmXLPWQNxCD8nEq
UAab5KMEGjgmQVHHJhGDFn58sbjXsNxPZzXZJFG2V7ta2CwPO7CYLgrt9AkrIlkc/wJXI2ALyqSj
DkJuW/kuWZ+lJNKU+oJyl1xHfya6OipdbwQipzFdEho8/os2w7rZNbBvdWL5FfA5qT3FZNwySYiv
ROKH4ivrqGq7ksT5sFMXyVL5GCkB03HAUbNZeOalwbllbiiiPZMSOjW8c2SkFO2B7ipecyb6SZl8
VOCJ3elswXvZNnCGRMT3556iIyuiupCVpW90Ke2gjg4QdJj7A59tcfKbGO16qQVngTKc5ty7UyK2
cNMrr6JecIj1jk7lLzDfiLhg0ASrp76jy6tBXtyFYm7LuaP8y1CbjHELS34RkGce72U4ukdn0SkX
f1JiNaOWIExpXsOH0L/oK2WGxM9Xh74gyjhmINURU0i1O8jdhidqH13khHuYGHJQe9Ah+yMeIQhQ
Wah1AC8fvfURz0yF6fkeKJFaskicAIaW8x4eRrmgJCw6bQt/S1hkm/2zS7bV3i8AsvDUV5A7bKU0
E5YA4N3XFxFK/92zXWWzhBl+b7rAfy/n3KoI+0rR98Fmez4HPZ4Xi0y5dAxGSDmmz0wlV7+HmwIe
+eajoPgA17delOYJBbTJEc50nPfS6/nquB+eGPE3fPP6JZSgaUDTvcr+bI604PJFnbqEM+9+1+QF
SRyXZhMzu8NPigzGTy0yjm0+qprZGOZICFvqy72YiCDgJzUE8jd2KPYtLFgduufo5Wwh3SPuAfSg
Zwb4ycfLWMKuo3c/8S6QA9PDoxj7OvxFKET4p6hnAh9G6uBDCYJ2r7TJHnOCbxlYNBLYs8tpA0Zk
z/ByTAFNvP/TA4pU3+6A1t8rFQaqbqQhwGPXrCpS/V+B8DEWg9ztLUCtCJxtMYos49rxy+qXmBlA
AfxT8pyR+B/KOeQWw1bWjrrI80DAY1QGOBP0PP5L1TolPDoikALtPXgR0Dx4CLv/oBpZHOfghLJV
Dvrlxelhzs+g6IFJmAz7fdNGsQRHsl8AqiCqAJAYqKTgLqtW4mwiKRLi+hzI2S0/FVSvVp1n6/Q1
SaeJRNbJ2sjC7PHE/dKnAP9SSDyzUnS51CAH0zvUeQd0n2/fBZEMpMO4P6uWqcUyPE9EZWrXNPCg
+2ETXRlfobT/Rx2OPOPa8Vd3lEoatBZJtODlojPS5yMlhyMZCtWu0kVIp6PcxP2bIjOTuMJNYCgU
iGBa07D6B/zXC9JHHXJnEp11DSh+SbH7QWr3ei17gofLtm0xPwmcpS0BBuhVvr0xvM8u71MD21uE
qkfQ7kXMkGtaN46M4XB3yR4Pf0nycvJdDpx/JR4q/Ms+V8jN0nAUyZLfWEJ2ZGPW1ArkJH7NyEeF
C7rnUnp0a/0W3bb6FJ31eiLRl7eQ5yx3TT9FPO6SOCdgv7e9gst3wSxLs2nW/lE9RRGgRfvOevyw
55A5PsGUd4kQKdjTirJH/aW6MWT7ZUW8jVpEqgW3neO9Y6gkLetykKZtG7F47x4qrOhvhACwpraE
uyjwCJnnzxIci4aDzjP3ZHTtuaT9ViaZvMH0sYBjaay61m5SnNBZ07NpPbCf73oQl6v56TUBLaic
NTqbBmKIuxmiyPUmuQvudB6XOmkpS54R563N+8OsofpmqqUo4gpTOh4pKac5JktApz/WzYj6DPIS
GCloIoUkAv6m51IoJOClwOvVipbJlUC/mIcXy6XtLCPmgFcdI7OxnWwUUGEuEuVITYdeLzdN+SWI
FwkiQszv5hmqT7kDOBEosUieR8K/kEzhGznRtM0xC1R72cAZ8sG7kjtG7vXyDxju3rHuVM59a7t+
U4G3cFtbxPBbIv6EnXDoQEIXvl8UMpd9a6FK+afjKs9zNs2O4DHNgxJ95EsX3siX/5rB3SGLjkVT
lAw87r7GVjvaVZy9/nUDUwvJN2zQnJoN4Da6wjn/tjKvbhNqfUHhcouyWOIEGFP3X0AOyLQdHOnQ
QhgFlJDTTxVKjAXpNN/6IbQEYXUS4vfYC/mVLdSAj/irmfSumfiHuy7aRLGsapFJN/YAmOfze5Q9
fZPlHMZtO7TFlJpfp14tBjan3OSAL2VuB6Nk5AKN8Q0oxkHTV64gdAPmJrRbvQQ1akYCZOgCjLnF
f/jLdN2bP+l8Ixr8Y9pJmp4fggSxkjeHRy5wVnNUYWFd+unRtnEMmXQ/MdshjGe/0eCkp6ytjZCx
jC043a7I1bHDTrAhjs7iAyV5P1M7iTekBSUFytLaqk0w5LwwmK4HyOUEsS6f098Zh8KExMScjmug
xrJUZDN4gPCUcg2IDJfudDtK/sPPtUq7AyJpRgTGQ+XjQEwpOcChN5A9t1at2+5sWyQxRfq2jpr+
mYQUGKQeicNcvoUvgqrdjGbNHTNbaXw16r3ieRQHkWjjwwGc5nI6C9/Bpdt3YXC9IgYm1FjwqQSP
QTlgfKBBETlV7ROI/1frJ6KF9t5h4ojliNS86Nrz1/PUKdNZAHakxjBg67QTHmyAl81CGI6/6sxQ
ys6iY1X7Ty0hgf2jigoYFHOFf7GGFGSFbaJ+jGAog0dJKtk2GDhCVvlErbGB83X2eRIg5VHWXI5o
F864JdYimCMSRxUY/rl8cRqdgvMp+mOLO1T5Z0BCo+N8w7+sRP5mT8SRBWX+losssJQrMF3F7rHg
SQ6S21yfNHbU98Digl0A3IXyiD5zTwyINa3iNM4Iiae+L5fAyeCVa3kG7geAJ7yzWTn7U/W9/wqr
gb9k57QRvoTp16DqGe15jR2kMJqHSQrw67vN6yKtiuVEA2g43DooUjO4QCd1AORvO4JtIU06zz3n
xBkCK9tQxSARDSMm3yyUu2TPWkH7SV6zpGJ66tZX1dVHkDoHEZdh5cnNycVTpwbX7Fc8Ng6tTDO0
jhitmiBV9PgtkPdrUNco4a1mWT7BvQhSU7+7HNgEanNFj698p19MrTlW87xp5kg6VnFEOAWa8n6u
vzutyaQROCaQJhe0GYeOejgiTReabJEbsCsoTWeO6SKyHrzLoAoqs81dwNclciuKnxw3aBXDC5os
Q2UomFaMm7NSePShnFFUrxa7c49AiFwYUS35vBSX76/aXBYsbl4u7nD6BJ/2N/4kFeIHEtSnE2eb
blPkA+zYVixLhgx+KD03biUTt9cYa3BpnOoo6C15EOT0kAxTv4eWOC5ybArrzM1QPxnqEljwJkf7
wTdQRLV7UvAvd9+am8P30B9Q3btSaSbrcmnGx8SFtoUBXA9W0xjdFhVuPojhiOvqBvxz/wHVpBir
crcQJQl9mqpWpFRtOMjqo49/lYVpfHol30mRI4NxOUNK7lXsnyZVLD3XEc9WUHQsns+P8zcp0aOf
kLky6BEfSOiqnAVdktNSzPJ06cxCOSXbvv9l1AaLDltEcnXIP8Z4dR2LYqx9rDF5tDbD/3xsxuKq
WCP/TJcLnxOsr99aOuHeeYWpNLgP92NQEQOuhvm5/tmcypvMsBFhH3U+P9YWVoDoBFNNXgZPU/ax
2LxypyFQPuntHrsdv6zoKHWeHbFfSTTGVjie8aTigZwcyhAByxAzfYcD2p+JJSEmwLLQZLQ5MDlx
QxA1XlIXA8r3GEovi+k7P/QFqd7uyHbT7CcQvS85zj7ZU7muP+qupXoyujBukyPdn2K7NoCP+r/f
Vv+/Wcyb+2xUs22klpsta7fL/igRexJlw7h0DTp7MH803MqDXE9s/0w2ASk0AH7HjUxOy46OnrT7
oyIjemFsGI4DVnF1nAhThgfA/dlzoAIQTwfoQ8CqFwgMKnVVQLdR+Y9xyQs1BoTZXQc29mb/dNp2
AVxavYbnSU7tocz9WqNWUvDrucwaeQk/EkVmNAYaoNHLTi3l+kN+ipv8Ic1WZ9gYBjUMltoumh/u
an6NKP2OZQ2XrLdaP/ZP7tFUv5n5GaOYmRDLI5XjRj+ZPD6MrCe8yIfLPxD9jiLGezcAu2tEica/
YXpKy1206UZATsOfdpdDRGqpmQcKxwjr/Ez+z32v34BgTroUBsSuDUmrmR+jwer1ArS5dGQqih0W
jxKT1gt+dOOgRgRZTsuLpCcd5mOeL0/PGPyUin8gihZpYXFqk7bsvzHIRa4jk6NM89aUn6Bj32os
aGzi+zRGdl+qQWI3F8CqNy2Bo5eX3/XzjoWOHwFGtsyjUC+y7upJgUWRfAiYPZC0rHrRrZyTrdRc
aZpoYoxMYbiUdPcEJf/37Kk0fPIvxIJOD16aiH97MD0ORT8NA3kD4IIMlyHF5IKT0rK+tL3OLrXh
vhR7genNYMN52OSCF390GwxQDqgUWDYMODJOVz4aICDIMtVQXeZYKI6eS6REawlBoQ1Hh3MJuNC0
WAUv/Bb0bIIobV14ehKsOi/QI6C74eShYBToHdKw0IjqV1WlbVUFrYxmid5YxeJ6xUNrDv/hqVXh
BeGAo8JeGNRxhhOhOWfoFU58V+0nDBjD12ZpkHJ56cV8zfuNAiNYTgYjjZQIYsy6Pm0fUWU7ltxR
mLYGYOvGKjMCUb3/1cYWV9z99hP9vH6wsZ2WSZqSTkw5W8EytB6nG5SgJJXYcrp7QI7rds72XUo+
e8iI1nSYA3OBhxSYLioYGszEuAYYfvEk3jXhOS2cPD2njz+G7JDbjsYXQQ/gazxShwMR18fzH8Ju
fXwYm9CwaqAN0cu6UdgJZFBVm74N8ckyRy3GNgMbeQkR9OliQJJy8jkqbFspvu10NzPuOOAHyg+A
HdSaYvXnodQg7ms4PxtPak1JXwAJdTgEfUEK9f0hx2GH0ZGwoq+e3NrV7pFec5RcUVyMnd3PxwuM
xrFYAc1TZ/pS4W3n5ZvR9qt8tpKjo79lTFkvFYPNDPxRwMSx8RSZ1I4EOysXp/0AWTe9B1CD+gon
eTN0Y71HBhx5esP8yy4zmfRjeQFHRpZcfvuCi3DZ+N+JyVlyV/2Ivvp09ySPr4oIvzmcvhYQvJXd
WVXMQBv9gw7evPWRC202uRxNWlnT3+vg1HS4tZIAZuTT6TdgmMymU4RxCIvuOEqch7eZtki6ZsTc
0P3BYkUvZvnPLaGd1ChKcllFcYjOI43eaNbAQ4+v5JVTCO/ADhHIikpevGxqLkwG9Ex51dUAnEsd
WzM1THLrY/JwU92ZIlYER2MWx3xOc9rZMQFku7AP5HWU0ra9tUcmN8AwvXi1BknwtbABI/rn1jZc
pLmm3w2nnm41nYZbdpilefdk7yEnCwoBZdjXp3pXdNIgubT39j4xJXpft9vBQY1aDxw87FvK12qZ
3/Wr1N448ER3VCoblJAaMRCQQV/MXJSAOBnpEOSKY/Ag94PLtWCJ3XubF2kfBV2gONYrpZPIpahA
ekaUWiO7/XKYUJ8r+8fQMude0DuiIq9Q87Rr3qcI5C8KhpPYMYEA1sVR/wbk5sORDciZ2s1HHq7m
etWawCYbnsLrdi3ufRQerFhppDvsY3kPgQG34Xka07oXT/c/aabfR5EqcMr4jcrjHiQKqtC8yK7f
oFpKkBERNO7cTK1MVDI8wMIPrp8/gvug7EfYf47NPQR6NbjBex6Wq4tI/Jr+HKMRsSluvvSI9DmG
OplDtxJ3j+c2NC7k9WLBL4ZCw4+id1WifsW1/wXFZzC4m9I45gZCH7IQYAkaKN3MlOsCBILhKq97
S/EpcbOvYt343GbAmoKDioqaTJCwynDAnQReGqnm6UO4qX3XbkylII+WiaHtVrm9i4uktUdi20C7
8FnPl3Sy3vLunuJdUJ31Cwe4Uws1IO+b47HD26tqzS3aKQ1SbmrMtE2Exd2eRa0IuiTs0GY40fcq
DJg9rAber3LeDXP1SqIYh2ho+JLC5FZ5PWjiDrZfYF2H3x4LGTwMtfX0Ti9/KGZx6lBRgSOSHqSY
vgg7O2Wh1q0atthrI4rdVeP2is5pflXOaUsXmOI2aex6dHwUolouciygV14wvS6laan20UfXsYsg
gZTPpOA+TG/WplsO8txkpuHvDmfs1bPx2aQIpugILM5dGZyJ7jGxev2nbM8zJOESmrBq3A43SJp/
dQgdB0PcaYgOOpi7+TzGp/6MlH4eet/+aiqjQ9hDF2FsTh5m6x/OHBzBOULj3H/jmlTdbKaGpa3I
V6OeXSLa0Ky4ykMjFED9eq8HpGFgyr4H1TnLPd1dZ6sS3GM6hNjstkRypwMIsxpF+24bWgsAtnhY
02ZbdLJ5Fe3/i2xd6FBBnJOWcVJ6C2D3xazE5zHYuOZNV27u//Cl5I+fDfwKRZXg0DGv4PKIHQhC
tUJ+3zraQS70CsCd8ZQNhgtSqRmPrszvZnGhgFf53ksV90ak8EaQrPa+ummMGrDjZB5C/BrBJb7J
bB5c4meHg96pa0/Amz/z64ZDwJ5QzXlUsGv0NghC4t/5cvx20D+ogSJjGLvYkTzEMVG210as31gf
n7VevGWsHAwjm872YEoQ28ZNjhldwUNX4OF3UVJwh1Lh/0pCwJak4UJ/cR36QjY1hPmrtHtCZTcn
SOnSaWuJyJ86JWqrbjaalYn+7T00U++o4fUjSgvbQZ5rt589VS83JDY3dAy5ztdmxYeQ+jEWPaCE
PF3mx0JNWtg1hy5tnyJdnY74u8RrcDR8QPCekdK+N+twiRr6reYAG27qfvay6RVQX75sns8OaPFq
z9LgDDgG2lqlWGX59DffDh39ZC7bfarVn7Fqvd+yDRbq/mEqYf047NeTMgBEKdCgZYlbrJiztjT+
c8jw9y8Mk2HC7VxDoPZxkxP3qFq69r8kTS9R7oegK9X29NkckE5MiteMC4mJJl2bBdAkCWlblADR
DMoqqsm4oo4Yhms1GjP5LhgYfTWoUhEM7s/HyDMzgCUeIRUMtM+TLPkIQgunhiS87vOXP5wOvIVk
8QzGxI0lGLCniyOuqMedTYeY25NO6VKl7/Nn5WOXx9euWCX0P8MEwNUjtkUejHoruUXdCpM1uEQE
mw0/ofU+mwqu3yHzhZXboBX3k3wmbTeWX5fLM/XPdk0FGbNTSi6CBsRXhHK8plSDVMHz4QFRdPxO
pjLOgBiFIp+HaNFbKeDOF0p7fCcDBvgtP7vUM9RpATkDVFtPaQfaviTuyb9x/OqUcouDmKlu0+8X
GJvRBXnUHoEeiLyMYK+lchb77MJwduYkqw4bPrS+Lw9/LK6GMURSLR57aMg8J3UXgLDjrwOndk1T
RDkNBgfIuCbgROtUcQsKY2NG0+veJ6azj9AcDb1vlTMToHPQ6z7qteX7QpXKvtBMDQAc0wvm9THe
Xr+c7WAkFy7KIeOKymTlPzNj45bRi/6QAJzZfzlmCSa7hQ8wAtPQeCfT5Q3X41Dwj8TNSOgG155j
qtHYTGFuCaOpl8b6EGcIAHhByEYDIad4abTXowKxQp8mkfIPqKb+JfyWOSG9Tno5zjtHGjqdw1ww
QbBfSWjCC2Ih/I3tD4pW/iRb3HTBZf9lyW0wc7UZh5R5jAJ/RhUozJosvL1bhR34/aYdC2ffw9Ar
69QHRz8ZrfIa4auuK7Ox/FZ0//GErCoYcTyO+bLor70gA5VwKGDYlRli8OySOI4WYU0HYKM7RvaS
Ts/A4iwMQltZbogSXOMS8IxlOgETHDcn/SCbGN/TBzSF5RD8ISiq8Iyzkjx7NyVd5XBVIdo0sKGB
HhVH+Dss8ZlSktlXpGY49ht90lIiaWqqwbz70lolvMvUfoZ9Tovl7sshPafwsnR9PNgCcmtE/W8k
a7KDx6dw0KPWIz/UIhBJLjjU+T0En4N78xfSpJypdBRnirzDQvD8+cpCCVrreSgrzEYzZqYUwLhH
rOUmeOTxgQiRDZOsLCjwsjLfvAe0dowBqbl4gXvbKN0VuexxNfl/rdFjD9GL/FgnazjfDhffRHS6
r9u9UAAI3xqLa0y6X+f2nuYAmVyCv8GiU+vCiM42Vr9DY8HsouzUh2bmVLV4gI3jT/O7VKTvCRRX
wNtn6wiTACjzz3EHp5xCdnA7psV7tKg7LI040+fkUibWB80+5u4QWYq1fp1wvWP5bSRwtKKfVQSJ
G02HDXJlEnQlztk3uM8O0CDAurThxhY9dxsw+96q3fPIk7oxjrnZRvLn0M26DjKtr33ZQSyd5BBQ
+NcZUPxh6rOPeXQ6slMIPLKNeH+azSWw3BZPZtZUPUThpm7uQWlqdiLKowLWEJbHjkl/GUwP+vfX
iRvefDqNOEaX7TZ1/zr4DMBtPHsE4ac4a5eJupoI0B7hcMgvJ878f0Wff5kj88XN6xJp7iCHhl2k
LNe6zekcVJMRoSOqV6hFq0+1h37YapAicmpO0ZsGp1HtfrMrW5rzsDKCYegz0F5IfRv4OTcab66D
jcd/z+k6wVBoTg8+MVmvi9lIp1IDPAiFxjj/b1iJy3jyrs16McT/0dJNi+aTFoP+IOutMfJN6+qr
pE9a9eghZjM3fKZ82YJxp2NTCRF1KSEnTPTzMYXk+bqpcLkhyUk4+j6uaINx9zC1F8ZYkE+eVCKY
J+PpHk5YM9JriFeyx9dLKEu+z26qdedOlt8Ay5PTuw5Xy+3nYZr/VWL22hgjzQEKth6qvmnRDwwO
gJB10SvH7BODdVGBHTzum7J8631pwIhf8rKto6PMtdnU+UsNFeqUKR2s53DiGlihhM3BGCwpKVXy
HR9AcpGcfPx2Jbz3xqGjOEUR+NpT2ZmjtjD5MxMh5ZBrUc6nf7qE8/lc+AEC5wB2MlrrN8xGM6lh
1mfuBBon+QEEydTSW2jxzJfNCT4mB+J3DPcQkW3KiBuqPNzyWO8M/RfVvy15nt3bpVgD0M7PApSM
Dt3gx4+IZNOOMIXMN5Fps0+0a+MwkpjP1F5r0zJx7UPYT90/UcNQ2VAM2ijSV5lBvM+gVlYsaPOx
bPb2iDfB9C+tpbiuASVbZCmFUa76A0zNvMusmpsxhhmP8Hl1XhY05QH51wijl0q/GjpBRNNqbNc1
PE+lDs9PNOzbUd9MJtd2OYlDJw3B3ESLDzHC9wcdzro3GIz6YavJbuz3VAfmCkEBQaf3Jms0iY1Y
6oGDzrMp8HiEuuwlGT4zDmSGxw0kp+2zD+tAvnMYToFz8Esz5dQF5WbOMuRn/Tl5xIhMh4gM6b59
ikQQI6253+FX+3t4FrPxSiEwrKIH6KqwR8iDmGznVh0hfeh1RlcqXFs7NG1ozdjZ4lq3tFp7Xlgy
boBpnNOa9QKOrb2C0HM2bRtOu7Fte1R+BKqyNfqwZVQCjuS/YHJI4RQF/LySt81WKRN9IfN8my60
Wy5tQar049M/4AjWSW+6uz/3KM0L/wpgqP3cnqr3RP8D8kTh7IHi3VfeSjKpBll9bdVJ8jaNJ5RC
llullnCL6ThP1XJPO8soLfHtNF5y9DSaSXU/hYw1LlKp8hzSuQBXS7gmGwyoFJVgqcUsoU4ybmy+
FqBb3QeY5aULs+3a4yrctb4uYPsNizyvO1xRlZDRceOJc81Lujke1cWjU3fRtBf7tDyAtNnpSUiS
yfXDzx65xOCv7zlgY9zuv9wyYnc4kY7M6Og6xjGh2Z4sIPbxqn6GNlZSNo2CmrlVJo/d1+0HiuIM
/2wJ+ZzOUE051aleOq8pjQQ3BP9xS0i7Zw5Nf6jCvf/1VmltCHa/ZfnfIAScTe0konZVWTjxv3Xo
PUJvTV5rSlGmIc+b0xYrwPcd5IRfyLZRZPvf9GIJWjfiFJ11+XxhHo0IftgbRh4De4mOvSle5uTG
CPdGt1fGhfnwunYIH5cZMS28Vb2SRPAE143V8wJIrQgqTOt4TKhK8jS65kj3jS/fvbN0qW3RyULs
2Z3eXPxBZM524mxb6sWZ+Z3VcuII9Ajd0aD8xsG9ghhugyFFitZP4HK6uVOExniEWwhTezG1oEFu
kMKGQmVby5SPaqHhLplKAFv6NU+OcEDTZJVgLKHb9X6uyw7f3BxhxKJ2MoPHXMy1UANHhglM4ais
KFcQZKsJV1CFCEUi1f75XZU/9aJYyhqJ1JwbiAOsxGgBoQhJJVdZJs0AtBWeQbmbjPEimCn0krNu
APE5lHQ+90b52Q21xBhvqllhtwY+Q6QB+o8chF/HeqTdegjd+r7+q6DAD1czjWqkLLlIvmo+Xs8a
LwrrHex2XcJ8nJa1PovgtKTBWAb4VTmw1RNIjt66viRcW5gtAheYZAt9ifCVP16bvad6pwUu3znQ
Zv/AvgAi2JMV8xT2NS/IEmUJR/ZTET9Swjn6Y8Z9rMcyp8SM/v/ayltNEt3Rftk1BmqKsQwLSJx2
wf0uvk/5fYlpbUrDKef6y5FGpBsxqBMb0USdX2bRrb0IoNlJVyvU/WVjJMFMXSbhYT9x9U1z8WvR
R9V3aOTI2XWYXqaWDglB2ieuB7w9OZNSuV8Ia0gxZMXK5Y8uOf8RdAhTfXB1W0QaLV0xliWNZKMr
Z6d8GuPQF1KslDvSPZaQ2d1nFHhUn5uOg71CRN9TC2ggS7J7R5s+8pcPJqRDw7DVh35jRHLzPPOo
KqZE2ScuhEcnKZksgMLNneN4VUoV/4h1S9QVidfSDjeUX+m1HnRgR+F2PzJPKDhVCSD1BS/+lA9k
NXM5c74wq2Gf+Ib2VK9sIHdqcgKMkRYnXuBFRKqztHIB280P7CsO1v/nq8vnU9eVOxnICmqmYnHd
eOw7jBwjaui6ANBTcMNHjJ4Xu7FN/VH11LuKGX57haOIDPeEMEnQWgFNjM3DBKKw00FOS/9Udsv6
vcq1k0DVhCWAsZZsAp6kWXO5Z12/ox5/uw0ircjBmhIn8dBk/qjEJZdLU5A5bWkGebJx+gYxcudv
1dhxENtkvOyQS8wP3FG8gY5adD78v6yBKya810NbusJguUnbWDxJAdbwT42P4LZmVeH4JpA96dkq
X0FyiBEuo0GClyvEW+KKeMsABDK1VyEiR+mzCSX3neczM1sHpmmR+ZwhOQSXqOZq670OHgCttbXf
Tut+1QGQjBBMaXCICh10mkeirJQPFaJDhmVhJc8UGIeQI3XVjH+GH/5ytK2n63DJuWhXMVMvW5Br
gMU1dD+tDUEexhxQvb4WbnzPtOO/9wD+aB/qR+P3DuFlBzaZzQIQIcmfotcj2mrg6c4LaOfsQnFm
uKgwD1Mm2Q7XsKKKz2tcyA0tl70/Buf4zyi+xvD6zUc503H4jUElL/AUmpIAz8jQgmDjQkf1otkh
4NFBabQTALqkAGADKJjbDrstNLab/6tZJX3PIFqnqanLaUmpBlUczZGg2upv2SETPaVF9T0VD6qZ
9kctpd8ciMj8MqF1tfb3ibOZ+jxtL1Mxtzf3LQBAASETomeWqI4lY/qn8whd5x3iOa3RZWBYSsuu
p7IopQI7PlmcYW4tC8izAAt8/jEcTXtBO/yrCrLY/WPthruK+8JzgPz4ntjJm6ht7MAtkwWPncz2
ugM8g2iSLCcYAWwul7kpfDTADzuIYN0egMR6p1zf2jQZhRFppn+olUjQEcSQzBBS5QU7TIDcXTMP
CyWyspBb0jgQDE67hd6e+uZoBk3po8Xe26Rsog1FF4uy+Euu15EfsIQdatv8uNHRlrUAn5g5K5Rn
IUNHZOIabf72coClwmwTbCtMpMPc+VTqp4Un30hZkzypkyTwpv47TKTsbjZiiDNEv5i/u+qYm3g3
1i0WXOy1ooi3adfPzVfoeeB3XywjXMK2TjTaaXH8CnEKsbp+6OcwUOPFvgqBp5ObSq+nPlh1USnK
TrQtHZVNcu3+eqgAjZCxEPVcCPU7I0slSGCXs0XEjVRuQayR+duZtCOVTgw6Cd7E9CIsB+VNfb1b
ls7AmAgpp6gyqdpTv8uFWJUwm3bLnVbxYMnebsf7Rj+lSEZ2LUoF1jEa3q0LVHVjJRIhdLx6OXB1
kwCDOR8jNVgcpz+ufVJJK8DB7RcbBqg7q+TtFdwZBgyTVF3Ggp/9pBoUj0Xt9F/cSMc0DyQsm2Zu
+tgXVO1ckt4av6MpJPInq85L5ABHtb7MParrbVvhaRSTMRnQFzLW1GFCyKTmDY+0PwuOwh0XgaBD
3s6GxxJXXq18hZz3U+QkDLpVEnwNA24yY7OSpIapmyHyhGNreHPvdzopLPlLxDFsRjJC8Xz5I/cl
Zgv9py0HG9SceHL1m2KE030RX2M+IImZYUfH3K6kxgyVUA1Zt35Mrue89SxTM1unZTWqeL2CutA3
XgNQx82+tPIjJUoMJjysoQ6qyABY5pBAItY1Cm6q1i3Q/YQNgV5iB0YJa92dQa3e8ZwBm5px3mM8
Mbyjk5VcLuDfozaAieDsp+lAcbsDg+R1c6srhQbSLh9wjITYB5IPZjrP+wI359IKDtUi5agJcVZ+
9HaBNaeWHc91hYa+kOMom1eOgHOcSeKkCTgckwvVpaRdnhAti3aklO/GB6k2D/RiSzzOpOnQHgRJ
9H8ANrki0WJlGCPJJEcBMHmoN4CjNb8obFfEjSlW/l3Sev9MmEw3mnfpdXoHw1rsH5OxcPs3KIGI
kf4LBHLXobwHcKFLi8cUj+B4mHTzSjggcOKXBCPlDIDHPdZJ35c2EU3S7a4pmyE2W07TqOgnHDgU
IpLf0Dvibtg/yk2sEztVZL3xhtyizQBOQWjcFJW2OS0rNFn3drXIRLS0D1l9dOsQ8ZaYXRmQ7DQ5
Uryado9NfCXf9AwRbmmU/Z8IsEGOkryG6KeaCwzfYKLAPzBGKVKXKOWK3c77EdUj+lsTWLzTGEwt
Lcz3IUpH4kZ2AuBrVTbY+mPtMaTE5LCoAujFZiZsN/qSvTBlVX1omxfO9YuHWIlPNwul9eIsCKoI
QNdpcb/1cG/BCJ5Ad2aFOR18sRxo6BAW6DDvTpbnBzP3ONcV+mpHDFOdIzCIfHR3pS38JdMRxi3/
2sIgVCW3YhVDP/lGh/FTi+KHBt7mmaPRWC6xpqnS2B4Yxo88DbQnnt0VYRDfxrf0CNqnX9HUliek
OtvrVIY3SPvfQnFCyA/ocIBU//GUI7OzjAH9RtS1B6dwARb2pFP+79IYxL+C5eexXL7wlxyZKt5Z
VGXsjlspUfNmmPKFj+Cbf1vPuFP75w3K8Z2N6yjJqNAx1Lutp3o2bGkh0/YTzCeHKam1UvusuFGD
t9F1pxIMuv7ZfmM5uApk60Z/6TridNnNfOgc2VouhYWoO0gaPmXVY3wh4qge+J1mvEQhHCYWuW4g
A6SUcNl8oJ7RBAHQBF+6vRT+aCijuKanpR4x9eBKSAxwE4lHac9T/P6YHJFttMvgpX1EGwU+VYFv
uk3JByIRb7jS42Q0tw7eJPaR1jahWAsUc3OmqJ/lNeYvffFgWPxd9gzH7snR/SDo/C1BVaqhzwie
UI8Kj8OZjTB+Nx4yCBQQkMUv2u3Y7yYf3iLQnpRbkX9xPNnarlSr+Ozfr9HTlLTXcUiIBYJSRS87
1qO8xrMm5i5lwTG1a6xqrZmYwiZr6tLrJnDGz4vUroSLPnX0l0dPinWH8n6joLpBylwCX15Lhcr6
IZNn4AgiLmRUNPg/mYkK+Rudc1Ed3u5ajy4wIONjJzsmuJiUTv8ZeMv/MZcI3IPt5LuOmyrU3S4p
8JgvgBvfvEuTxjRkYtYdMtxy1tX/POjv+7Um3/bC2liNxqCY/CEyrm+x7c8yjuFytwNbdJV6RgQw
76w0cUkn46HBIXD/BmTKIYk2IIP2aouGTdloVyQ+FmMj5xsAsUfhk6GeUYAm0G9ltsJ/WjEeDIN/
zLRNtn35kk+KUl9InxmvrVMiS6DWV55z5uv7vJ37hXl+YDDy22vxCX5BAAX7lyc474djKI5IokcS
TymUVKIv8zBMQycX6xpe+Y90iOzahJphGATdNYwonPiSveABzaouZFwyrBOYkaZx4EmBTKMMcBn6
uj3gwd8YaHumOKR5tsoaBjEWKesSnPN7LnczbIa9cE5rWh5A5a5BqxHyap8gvphquSukS/x1rtv4
923Q3VqwmTye6HUUbkSWFpWX7aN8u+598TW0FyYxFNiK8V70IOM3dawKihzPrnBgAvWJ2KMOHg9a
zpeDiKdScXlllH2zXYMcVWF3h6Q2hliIHN2cUeshPmHhDDtT038O+sRwnxtqOfynx1q/snVRIjYZ
HB7oDCCJwaij0nY5g6f2a5yoaczTvLITL8Pk0AUzT53MKDmNjR0wWUHi5zXOMuVZSffwvxEEj8dL
rTIvo1OOvpWAXz2Zs+m+CtTBk7TdN9BM65g4TEcoh6WHPE/UsUUF6bPfkbP2rOrzjHJBivnbSPac
krb1lNOjdfpdQuW3I8rQTxhDo0qdkdkoKZgXmmj5f9ZdsS12PkNl10jnMnriHYdLPWDN9XkXbTAK
lgwNcBpogGvG4kCVUDQc6TZG95dq/qcJO/i3b43AXkuQsgirn2qBrvC3DDC88vUZIaUIb9LVGNW5
UUU0iTQY79poIAXfgIjk8VftRgisxPShlaMpGWol1Jv4ymaAIma0gbp3MPmvACQy6o+Xa0BTVqmo
0Zxs63Hih8U7DCxLUK9jYVjLW1EEQHXHKv/Xi5IsV7bugrg1ByszZds3M+cbDqkQhP3bDaYq2dGD
2M2ZqPHeZ9vKEeNgc19AkJPz8TXbnVquxHxsyrqpN5Yc02VvEeMMwNG2fHVp475xMLb42vEZ1pJc
ncmOL+F7NyQKNJlcMqKY/pXfXxJPag/KWlK1ZqMtEp4yc6seY6pa9MD0sZ/Rt6m/OOShO168or21
bgpC++zySbS90akXCuiBhfgjFRapjhBu0DybGmHeuAkI/cC0JNdlZiDNYzrXl1daDkzevRbbjRJj
VD9Cb8625PpJZWpJMnyjLkwKL55IdxphUBDMhO07tGRBtKoPojY1LSJ6G+K0nJgrQiJro3ca9Mab
D9mZbKjk4T97ojsMR07MSIRt+27AomSplBscGn4G4ED0a3ufTGG0ST7dD7SAvY0MbXwoWxjXpibN
9E71/GSal74cwNe5xCKQy2k9viQ/kT9V+RmdNonFzyHmSsjLvcLDGm3CN4wz9PkEyEwdQhe0a21f
4SO+JCscPQ4RowyXOb2wi7s1P9HV4uKcBSkxsrvY9ziXxHBwf3MMqIo0UokDA+I/s8iMn2UNHUIp
p9oXMYNQAHrQhym1BtSwPx4rdgCh978hqpZEdLARSUwDqlErbii3ISO5REowCY1aDqLwUCfnc9zV
quL5IqfiR/DHYJc3hSe7OY0UZg/YnklPSBOhr6bmKcSFoLDMVgNwuv3AtFvCwdcOROMebR7AnKRr
g0W2+y3bV1gIl9RsZnG6Qd99s2JCH7x0xC8TL4H4rQhd8Xk0mEaSJvhtN2tmWckdaw90Ow6U5x9f
qHPqmAigiki7P4kcpB6PUJ00dUwnoLwFQS+de011Szj8RrjuGiskiSzzEafPj+84+TrF3npjK0jW
76y+ItOvt24y6pNn7NKy54ce4Ss4v3mLnQxbgwBAwVXg0pjqCy2o4ePk5cxhEO0GGSL6IA1fZbYE
g0+MJLp9bhRJ7Ktr8W1On4PrX008TWf1uvFWiL3BPMJVCUab8rMWj9qJRuGAcupkB/sG4eUUdJNm
DxiRSK5omhSVdKRAnJKQfagVrYHnwpslgZRg4L9liO3UoNHr4RzMAda8wgUVgsX4fzsLYDNxmc62
CS0O36OI9wWGk/Iw3oaqEiHBM8685pzkFdrWL6BnTd5WC1TRZJbZ5bf+cMO6M1TraqBmgd6acPNA
sh1PiOlzDJlgwpwcvLdz2G+4E0CgbQJ9YOfmdyz5L490eT3mPv/YcOI3TBz3WlGSQu0l3p1z/jm1
B5RHnpvhQzWbZGcl5Fq6Y1lVXNGzT12k2NGMjJ2YAviDhh+bZxxMzhoQVFfOAHXjW3BCN4v8cf4c
DBk8RkvrvfSF0nJfwF3r9zyumJf0MI1NL5NPfoPZRuPCANppo6Ai8MAgpn79uqqdboQLeSKkVX6A
7t2KMjLmDEw41SbWFbJF5TSl/fTAOUuVCXbBIpl4e0u4T7QUTpAIYZ5OLNgDEn2KsH5j+1UD1RR4
H7OoDjktPx4CJnFp1P49rFjUF1mGwCdv+J6v8joerES+dJvFklvHP4vH/wKcrFwPuOjmwxG/vg4e
y3hfTpXlO3DAy8IhTOxmo0Z03uTTkSCCJdFg0vMI9EUxX0EBxCWvVYeLxx+UL8aOgnIKPdktxgyY
4kUlMlrmoFdDoBtQxNFuR+k+g0GROKV1L2Gh1qOe0DDlWGY9ICfBoiqbWCeKhZVYT3QavgpWqG4r
lG5vWr3WrcJFiswH1G5Ji38SD8q4qMYQGJDW/ZtC8KgvVk6/MC5sw4Ygez1wYIQmWneoZWfZ23us
lUH9Go1h6Mk0VUm8eIrqg3YNzo+i3/M3a/p5wKlHLwV9fBOFurLw837PGQURJ/xs3XG8KqVnSzPg
RpRbrOL+mSb3E5hYF+4Aqw/ZPQy9kmud1tUXLYo8Y4jT9gfbwyKlFCLbXbCfmL2+E5kyGX42NGfO
IZFhPDFeT43YXc4VM6b6cn2/PryaaBcQqTcQYWsv/92LDybXw2voHXsdSleTPfceuksHGqqATWNd
Cv5qeAlVbJJoI8W/oFwz+2w9L6SsqfvCO331Pa5zZZGQYf9/88tEzS5Vz46+eW+O26qdy9ydV+WS
04YVfhv5RisAvS/BVWqLve8ppc3Znqu0jC6vaGrmKT658zvPm+r98J2uU7scMB1hFIiRPDgHg1+4
eDpV+9GRFCsz5ZwaJBkwNualCY+t4LVcj8EzHgPZyyp6R6uEiLGBe4QX+bpQ8ygUT2iJsTwwsm5Y
31k9GmjjyrWL9DmB+DiQPf0u7J5z7dECSs5a4HOeZYQuxeZYEto7FtioKbsE2Tvsw5AAYQZLmLXQ
m5aOwr2WiY4/dOkMDj7OlLUogv6MUBL1JjTkttkUQZImY3R2jhP8ktp2cg+pA29OaoiqayHD1cof
Hjo+XxBxk8n4SWqXp+8l/1IX0++h4dPDA3pgq14qFWE3O+pQgyFuxd/BO4ifgCH9ueLRawZCe/5T
STFMGs1oxxuiSD6IOFUyvhGoukkrFDh3c2ICkHPPnczer5czM4bieK8wTKwoty1X+az0sxRTt4/3
mj8nclUDbYT9wCoyHQ5twMgMq8IPMLNMmdQTuQrw3NaPe0LJGjCMWFJvEFcleylgiu/F3OSlgnAb
zzpJ6EdXgm7e3slAENZLBn5So0NwtYqcie7hezyNEVLCsWoeOBuwmEcERl8iYZJaGiRhV20Xopdx
ivc5fAf6c0o+esoUmcjpbICHsX3UgSlA9qvWAYVgghLcQhDLG7Yez0w5PzlTroPITGihABZV3VOY
TyFLbxRs46xLBgYTgb8+CC4EYfLRNlSMgtTsSMVgSbFqch4TqN6yToP0Azefngw5Q0ly4HgXvCea
E6omsq6rYUR3rt7ZGbnktzyfWSAjUlS1N6sxYhftnG/4TPdoc2dhqN5qF5IrTENHvn1LqFSoA2xL
C383HmoXQMb2HDDgLPmmu1I6YCaZJe+YfQcOnJ7XTHzHDlgnxfmQ+6gvO7LDYSj/80zqStqm5QBp
68GrpbO8ma1gHfOJpubcsJggPbiiSpIJcKBUkrLzRiA1X4/idOfwnB0Q75NrR80ugC/nfddQULol
2cOBiPF8y6hVAIsFLpplqwjVD0DD/a7JGndHRA8iR7aXDci/6m53gOpb6xKaeEDsRzxyIq0EPlin
5Bxv0uGv0LGf+AdIfnu6Ry5P+UOV8BzDd3NdCPqH/qVYu/yGmrK5KPg6rg6g/VkBRvpo1Oc3dnMV
uniZLCS2bnDI4TJKnNaroPG/+X0D7GlbQA4tS8/y8BZmSRaGrx0uJmdpU6ruSo+sQtBovKl7N49w
eJ7JLcjtMetgV88e8LR0V7C7KkJMdqhv1J/tGWqwJ2vhhX+Gc5DlNoAG3Ts97L8rE3X3Max/kUHr
bJOBeDNc+DCwa4VI7RREkkFkJ1wNN9C012DkIAc0LnI9sLXQPNNU9B+CjcEH0esCHFsUqp9L1a6A
qdwUSma0Hv+w8NMLM7BGcvBxwavGb46+l4ZSUWcu7k79+W4UbUOh98NbnXfy867ZnbqcmwdWHKG0
DWEsjOf9MuiAsr0BaeZ1WIh/8ulfqf34zu+GgZbWbBa6CTKQ9PZTs1OOQjrB2+RtQy0g7x/VyikC
Ao33GAzh0l0CC/aUBAS/d0b317sns+q/9fjYT6JxnrEyjr8KdBrTPUdH9UBxYDvkuotMZNSotcci
BEMIAr6teNW3FvAEqwGbgQD0Ccl14tyxDtb7ri+srR/FWc0r+VwmYEWoIVnT0XVHKZPtSjmJsIog
8x4JR7Eyb2JFNkmNB7bPGof2BlHvGEHLROfazsK5Rwt6BHNOEj4jBoKT2TX5L9LvWx9RBbglG4XJ
jZELmXLEQrt0TbraeWTDxCeTyisZofd1amRmSCEYgTKlOQJYrChdD3unu/SnCl8axX4secSgUhwY
cHaV1sCt9GpmBhFHdu0iCkWNerR72ulomZydTTnGhZKEN6GxGidQRHyjNnD/LSCdcO1kjhX4zufe
mWj3bv8ffq5wNKKdG0jVQF4nzh12oSiWZyyUSgrzZaSgX6xrqOPw9GrR/psQmOyTDUeDg7NkjKR0
MpZXn1aOCQMoQFq2NZf4b9ZD17faY9bc5wOgoPOuJ7tZgmLUmY7Hn+Qw26qdBPM7BCTeOyw3FM+7
rnmqmERwRyCnz9QzO9pOApobQw000fV871pIyJM/Q9rfPC+Ok75kYJTJ0XTmYCu4iVFcx7LYxMFI
57rlzOFNLAFHVIDOOyK35iAHXSJRfCUWn3Idp4NM/0JF53kQmheIQ5yLFuqXWWvLpOjiu5lzTEUi
qJ1aRSQYRWkepX0g/2ns44L1x4kz6Xk4AMLQnrf/hIJmrWDvw2yNFiDgxambR6VwpcW5yRT+KklY
omdCGpwqMJAZ5+90oGdDRnOrZ6VTNTM64YsCCDmMI0Bp6CXUvrZ1fBcNb3Y1SbMrqSYPH9WwxYR5
sfAT+y466bcDygZB3wYT7tk1Et5TaHmJwaJtzsv1rUzYLo8S9Y4D0Zc/O9nDZQMNpVNWZTiSRZft
DUc4Rop8jtU3+GQ6/vtupgXTQ4NSV09rvi5mvLefcdTPu8LenNeZuCHyWfHnJEN4lsU+7Zb+4niF
mlEBtVLqkU0pSd20w0DhVhnLR0fScNu2JnRUVKII55r/JdUlnCZFBQQAgvF5+Oq+mNfR/sLrNvOV
EwrhJ5cSu1PrQA+4/R95MggnBSxTYn1toQssKNKu/ut/QoxZWH+k4dBeH/4t9EgLjOdsfp6PiOGL
9ILiSDZSce+LkwpshErq8fga6UkTiqc7Q96zEg1OYfAqpGQaDPofdOrcvx1SfT2rOdS4H2i1JULl
tBbc+nmarzGNXOgaGqyGwcjbJh0/rjWmhw9RhFDQHODzl7Aq5Hz8G/Gq+K0yLgHT+1+oPGJLNIxv
8551n6FVAT1RTn0TL1zoG8787qhH9HHEeM92uEgVlfZTiYxqO0LcA85613467Y3ApVXGuQbdnTvG
nYOACRBBSrLbqaBdTi0ZtwyZfXXhdRStN70cGq1+HTd2vlxzcguD6QuBttdSg/yFf95dLhbNlltF
JUB6IeBoi5sxgiImkik2fzjz8nXxBtKY4sp0ttNfsn0s0iq+278z6/tJl6sJoqofQx7cMyr14+76
/BWdV1Pa2WUjs485BZLFw/wFaV2bGJ0/YZhNlNp1PSDqNpyGONblQcimKEhwOHrho21mEBbXD2ol
y81M99+hZN2GsUBG01FVUqjn14DNWG8I0YDjyHtwe1N2pJ3g/VLoRJ1NMAhQj6aUc3AljYuQTl10
iyLhB0Of50dlLp/YOenGnYNXD6LX8GhapSnLbb9lOmDacWcC0rLPGiYICchG6KAVCQSVhBy4tDpx
wBWOCdu5MOSp1+HGCK4pfVUROMcqXNaWp3xJzZ6jyUHkSifkI9QPqcefp0Z9xrZlVDNaUp5pwwj7
p+qURkhnYRXWraWAARRar5h0hAgkKMQGCuxgzRNkxLPjpjtiPPzp6NALYBrq+PfpLNqHnZg3AHZ7
utCgtyXfnxC3efen+Bi4brSbpptMnpuny97IO1SptsXVDNRThjeF6OBRri3+23ySuPvkkRgsDqlU
QD2Lofoq9cFlqis6o0sdsFyokXeI/tdoXEAANhvnmdZV3FX1ve7lJmhVby8LssnZruTmk/5EOINn
Zbyfp/G54F3w4d4gmWdgu7s59R4U0khIEwJK3Lh2TRfRL+HYmBkWmjHGHhA4vf2tuaD9tP26YCu+
auqxgk3lY3k7SqDNEfzc7uBwOu8SnU0s4xj38Hy7NucMbdqwlvq7c122290dAL8Al2pHkUqruhiI
DPT5CEUJDdNyLylHm+TyRLRPN/cSZuMSVSw5iQ94YrrKJndd4ayAsiZxAoFZ3s21NorohZJwWJi6
yC3nRhgDQndBj+wSacanBnj8BMW11KMTefxUG5YYUNZbltfUxt2Nx+gmmt3+zFEZEN10jk2ZClnr
ywVrRNbbyWZ2dpouG2PN5ouyObzctBSBOeZCjlsLtSR0lLWC7C7xRE2HJWfeRpPLSCNSnzpMHD4q
mI+X4vIOBWDK/eMauixX+LZSkW14z/mWzUgNlJ8Xx1qUtRfGWUSw3xwWVFQ+jqXnRW6Ssrext51G
mEsmvi3sYPdD9qitzEf0bDC7Ife9o0WrXPmBKQaxT+dzM5D6COD4yp6BqojcUOv1s8S6B9wvNAar
Eo/EdvUWBmfEID8xXwbBY6TATTMWjgGTH1As8nmpWRwWFN7LeiqPJBfiv9RJW6GtPmsJxhJjPPp1
/OYWb+pubAH9dWjOzurfncSZHXq+x23PSEkxfsgaD5Yw0qWAyEC6nQcHWV9aKS7EuSLTKD4pcZEK
2X6ZSI1YxvyO6Vf/jw+L6AlLFKDNVWMM5gKH24SCHcqRrvcSQnQbL3Ep/8Xsc8FOHXkJkGG1ZdBU
dP4wGZ2wFLbz25ciK+BEao39dNyXIfiRH3kukH9QW+lOZl3yzDE282bvER6Tooq8pJjT1JZApCwT
QhOnqWtG8d3bYwuJ9LMDSEAvGpUbXSVuFkQGYPJvLMkRz9PxAwgUgoR+NeBRU2VxzgRsmJLAWAQs
0yN5J7+NDLz/42hB2Ohg9EmqYdmSU2eJ0rJiETZWZHxe90fUvBexYS1KGV8GWUyLRHJhMoeR7G5r
uWt1DSBY2WSEWqyCq7mYfCdMPVOC3rwwLg5tKHfKK6oqF3MJLU2pLWeFKG8ez/JAAi53rZ/Yw5WA
/+fDFfwY0mufL61ixB9ySOuUtCcCnu8Jcsw92NuMgRhiuAaVvR1KOQC0VLxT8228FTYXFIl5EuND
Ea6MCGRUz6ZVMsW+xJGHurtWbWlVBYPgQ+U3EqXbSaZnurMcXNtbtXtqIn3piSNtsHOtZgY5hUxV
PtEjnJMebehVnS1w0ynsABns74k/eNM6WOWZvJeVEQR/cMVCqIo0HkJMDao0CkQhbM37Z5Rn7mpw
fWI5++B5UQj1Wvu/n59mWcqX1ys0qeYsHBwQyleWJdo791xpUMRmhb4wq4UXWulxwl0lJBsqHhmj
S8mAzIfp3xgN3/7mhck+Hwvgeq1I0LkQLiuNcTpjHgJ788lj0ljTiqyJB63nffXDdAKyRwXSAMfm
aqqMviXY1EVa0c618mnWUW723qFJiXRGKQKcFBuQVfTKiB3JsN7hHBQ4YWX7fBPugbHFgtsVJcAf
c6XoRuYVDRYf6MwyU5Z5XGCmgol7Nqwnhlu4SOyuuaNFWvCFsa56ZztAe5Jb1AUFDOI41KWLi+hd
XZWOaSowFh0UUuuqCTWrl5PYMLY20tyXu2WJLfXlMK67QwGCz4WHSAvzT4hCf+EqjhF4Q6QmhFPz
UR6H1MKD7vLFVxTlUNUiwH//1xuc2BlY6P5I5NTwwrd3A5+AyeJpteBiyKTBgiZ7TzP67OFDF+uU
kIC5Re8cTuFuBb3SOs1Y0xtnIWqei9HtsXITQoP6dZxZf4NoN8Jt9yud4tOQ81In8rST1bFz2jxa
bZI5T5K6tIbL/VDGi+Yvx4HY8omObJGJcnB/jPIX8O0YgxNGPzDPx+e+il27V93wwKdzni5ywj8v
bLAW2+ZdCngRQmN9x6ptMVjrOF//8Uvr0QUqAy2+3dr6lATS8n1sodJRGUFhOb2I7B6oMkRtmA43
MoqF7UtoOTwrupojIDPnx2aWyWhRbOztuXH16vUg2zTFOYnXtuRiVPfx0XbrpvSzk17AfXtQcGaf
/JYkmYJJoMG0aMNSmG3jv2B4VkyYT6eFOTjpKa/ffDLIrQvc1zouvAJJTlRCPJS98IL+nZXLdsnX
L67aJJZB1SWDe7PNt9m6uSvdnbLB9EWImO/v3ibJ203d49GBoWZ/wNzYWU99JlUYkLgimvr1LUn5
7GOig9HdEOaSIUz3rGGPtfKLgFHrkZZFoNuwjTVEpVEol98LkDTNTH5UYwDtr2wYc3HE3iRTcJZw
lAV/3hc0zqJL6y9D4hgm6VRYdH/5iv0rivpokg0ZR6GmDHAt9AD2hwziHOoOtfBQswqa5PACY0zV
3s3jeHCi4F1SaIKCYyNT3as8GeynDV8SVs33IYjsw31okoXY56/k3GbzGcNckIBbbzJgkVVWfI57
/P+KbDFZwkf5BmuL1uHZjMb902P749tR7w5Uv9UB199f+RnyWtC5M60xb7KqM5kTnJK/jb4ocNMG
5v8lSUOBmJnu7XE3h8z6DDrI1Hlpq0BnOhejG/PmuZZo09PcAAbYdjHX+fUlyKsj7kGuhwDlbbVU
OUvxiLJJ5bPQb7VmadEx8vomwY0qgtFNwcCmR15xAMhYGWKxgplYAetED/XQB0+g8tG/SIzUpqeT
xP1tlSWdk0n3n5qVN7coytQIAEQK/UQDoIwEPzwftTqISSp7Q2Kqv3bHnE7ihR7sZo/DWQ6dVC8Q
O3k4y2uhyR807rgRmC3+TFTbp+cbRSik0+YWIbzO/0SeKLTanbAb+LhS+hVovaug2FM9KBlFswnQ
QXJI+Vw/rHNEhc12X4oz9kE/RMnjzXvo7kkiGdPsCiJeQWNcEcrh8LYAog9fNnpf/wtReLBHAw8o
EBDcvdwKaGnYq6LDPe7A8FyIVQW0UvWjlLQogI10S0HAmtEayaBs1QqqCSJjTCGqR0u9+TC9aMOQ
veqXq6svlh1ORp6bhDUnhAAeHRMtIdI8VvilRjxkNFPCRpY+YLQLyuZtiVY6+U9yedDi9tNIu5Mu
23qjL5RGQUmiNVNDd9lrU00PMn60RxrvJ5jKxT/KDd7BbYdM0hSnh9BW1+gpwcPrXgF2UznVqLsv
BQbhOq6HgUcdlJgcKszielQmMFUeY9JR8kRB56E0lbUAwU/VKY0iFNqW9tfEsIigIe49nWKpPWh0
yDnXNf/xKoQYeXwnfMYOwUG3WPAwNrQjWoxlqkvVnBBOV4w6P3Uq4cA5eMDKs0c8PSA1hMhKdEYG
mE1m/ePiSuQtshSvBaaiWMXoLM1LlWSBFNxY54aCA0L0xwNsEweXPiZ66mAEONO27sKUTT19jdRo
kHLnTe+WyvDqyBwgKW15952Va8b3hLf7jK5cB2Q0EZPI8KPHRVEtHS5nJh/8i7JQQGooFyzTbRgn
6EPXUmBXeh0rEUN1Qg3h8Kv/3Jiyfou0Jd76ZSpxGkfASjLp8PELQDsiNM83+6laiWP9mVH3SVLw
34qBl+EIwdQJ+vIaYaoVpUFsUrnIcM+UIMd1YToa5SYTrAwFJLIUKNuQc9y3H2YTfMabJYqB/xbz
g47/32Yw/n4KzAHdebQT4vN1uaC5DO/oChWnlAeC34Z/LzJS67gNCV+yeW3pk9cObZishe+oBRW4
eUh9secnw/w8iqVcWwHJI9bWjP0Abk/FC7yu+s4orwhP+FWU61Vb+eEbkVDWTETH8bw+a9hhYRdr
NM/3qw3IopT3EglcR6b0bq2CjAOcNPe5Wlb6xZ8w3nqHIGzGk+iWl/skQPfHtRNnCcrNXQDOAALL
LROx7XLalwMNc9Zx29aoBBnRtnskhgJ/+6/0PPSBAHxbvud8k1KtIG36QnmQXRYtUrkjQ68cjzP6
AB5O24y6yXcMUQZapiDZ7U5jnpMaED9coCnX4AhUnFGwETOrr3wlzXWdfaBjUvgRJlE63QcBOxwS
5qrdc+N7sPXJ/J2W29TRsSLP5xPFwaQlsq2NYwf+usZCUU28SbkaU5j9Vs64PQTPo8iHy3Mdostb
Sw/acRU6UWUY8rCQh/+33nRZVEZzc1PkctDqnj+1gtJAMaHPt9xDGy4QDTM1pMGBgsLhTHMp0pMJ
qnaxGuKoJWyXsmiuijqaZJJYok6HoxI0UgvV1PjOjHEHnJK7qEI7ZYO8te0Qwk6t6HcseJz5Qt+d
7cttkS30uMYXJKhuBOGSrUk9do+4s4yDqT72Qm3x97V9EgUTVjZ+GpcSE/tsfYMKzvDZf3Z0r8bN
Qb9qPdDYKiOKYdTCrO2Yw/MuQ8D0VoHaEJIG7DKHF5FBHYNe07ptZmOGhPKW0Bo/4PbgiF1DaUTM
gql4bFOKZnfHOwavaqDW2B+y1ZNpeY74Cgy6IbgVw2PwPkkV/z1QV2iIOoBM3buTYfN8kxTgK0tc
95bluU+E+t/npOEYdafY7KjRT6y5H2NJLoCFEGEd0rDPpmFARz5Tdw7L6yxBkbM1LIi0ren9wZGJ
0oUQXELHc7mcneCUR96gqTP6AJo4pSqnYPYK2VkQnCJ0ATaVMsvrRMF5bDwZB1nZC1shh9ZnIfig
K4wVg7PLB4MSiDi8Dg36ckzSaJKBw09F2Bzo++8bWWN2rFGHuOUNTZYZNFq3lXC40IaLps6XVt9A
0PqMd6LtaHkNbP0zPF0hCayGDqlZ5YOtkkxwfVXmBn8//Q61Xhzbx3FN/dZaymeMRb2LFas86kLo
I2cSDSdIB7LcHVBaCFczkxpcziwcSBRhcLIdfmBTnTVrMCptz80fV3vsTynEOSftBp2JwveLxqhh
zQnUdsOq0TNGSG6H6m5ilkXKvc2znylB4kyRpITChTrlr/NcQTzDnw0BjD90nsbvBvgCDvEe92As
CPhed+UmSAMZmM29RklKYlFz7e3F0QxzvXENQnH/EBN9qE2oHMYTpA1UJ5NsMQP3YKIH7qqT9vDL
8yGAZ+Ux86uulA4+MM0JOGu5gPbJahF8yJDSLNBWGoW9+XwlYOmOPi7qDCUAko8Z12PTIAfoNIxi
aTRQwCD1GCsJzCW0DIk6B1zR1RfVlvEx+110ORhiuqpW1atAUD0lifkc5IMgyi8+xVcKwvJH75xG
1FQNv0vIYowMvmTdOQ6T6d/krgdiBzP+THI+KAFVC1yCJSQHlnP/ZTl9YxVzzFMmFKQAaZRkjNUZ
ZrEp5bAWY6ZgNzg10s5x5xvG7T11GKZyfZ+qU3yFfoJKCY9wHzQPilEj+8IfLw4LnuXY40f+y+h2
vdHkF0qyDfEAxsobepHzVsBJfq5xkwHbl2PskAYKCS9yR3qGGc7wFyxVYWJLB0Ip7rd9kLxusVsS
2fESyMh/8IBgdG9Sb674D/XF79Dob5yUUMLqxg3npXfJB54lXBrgDmFnEjbR6rFh3wWdWtpRH/X9
KJ025Bnd2N7ajyMMQ+NH1tYzmdauef2ZjR8x1sJowJmRkrZLicauxzWsScynRtlQroZa6fVbNHLW
133C2WiR1b7Vo8qmluXXXHdaCC1DyAJi2chDvubkzZTFIz6f5DaB0pH6KnGAYn1o+NjULhcZxHVc
nXPGlyU64Z+7FUE/ww3W+bLkJtSqawMXuDgAZbnrGHqgDkxSA7+ThXZrICNcVTxSfFjWL5RN9FvM
ZqBHX/fDzsbmFNC+yO2Q7EmNiymbr3kGaIlDUTMs+LXoTd9fwmT5r/zsmdLlOd5xyl2G6pOfEdDB
zt3bndxlbnCk4WpUdZfxdpONzv6SGLSUUXaOrRGg1fqn1SyAI68jRJi/CegvWa9b4iuqt1eC7wiK
pEdfDJDm6Miq4ZxyJDxFSL/RwIbXPYVHDh/OgdLj1S5yNrq2t45Prpl1mKUYhEVC/NGYxIyX4ZPN
y89M3fZfX+n+4/ncdH9GxpPyUcyRuShbvClT4iEspaovuRtPPlF5OuxIHR8Kqj9bWbFzJeYNm4N2
bxHklkm95eKwV102+t6wgx8NsbRwokRg7Pa5mGd3+qSTX7IjiN72UeRejaRIs+dfoHcpoYRqqqXY
0wSRRHhlqXqVZkT5eOETWn/65/NZgmuVoUVqoaX3DKXSmGfnLTb7Xxnd9+uTJI0z+AiSfHR1ZHkP
PVTumJNVr8M/lbI3CW3zkHCzDPq9Gm4wJ7FY78hvua7iyqgLXdREIe30j6DRou2o8YPbEv/rzAM9
RYO8ehDGKXTiuEfRrUWazFpBsqie1vnFGPIqxLtq5UGZxsTVeZjaMim/zlQZJtuxfWzzFFO6luDT
ihZcK/Q/y3wTFmMfGTBKvaEtxOmtspDY0esxl1gfft4ir2CDJS7iV2mGkGx/UKh2C0mvwf37AjzX
LkE49rISCMT6/Jpq5Sv+8R9Fm9i7SnDI+4cPvuo7sbMyTmIVLDDro0ElL+8YrEhYi1EpEyV1St/3
aoWloZbvYz9TPcGgplYA8pElHfuLZG21+CZUr8Ew5H7+2+arUIs1NbdS5oc2u9iZSDeltrdKIDRD
dHBjh+ftKHXQTCB1NRZpbHVtzw/xTAKtenxQHXceXZYqQgD1G+hEntLyhu8YeBzxaE0Eq7LTa9+T
ZlH1Lary4yaTV3MsB6miXQhQuvQN2w7hjF4d8z8CBb1Eh99ml7+/3Uk6rD/AkL9aIDnVtvtK3oB+
U791OvyuflLGclTbER27w4DQJPBwnxrnR911eOFb8KfeeMckgwOLTpProet2NWU8kyrbvn15XsST
zz1i40doGNv4weh+9RIaoVUv+YPkgXc+jjXX+uJuAVWlVNffs70dUwEyqf3nxEYrbuDmD/Ot0ZSH
5CAQSh/WIUNIRnmwb7G6c4bifoFuXXGthh4VTYFQoF6dG9hodOEP8exdwAcVKw7PuJfi/BufD5Sx
UGxDuiEKHqaL12ZPVwgmaQiH1BL7j3farxJCPP2T6qAcy8AolwYJw9LocT2HxgNQUzHAYP255G+A
SzFvmBEdC7yxk+hhGhvPFaNKg477l+8v+h+dX6uVRNu1XWgsHxC5XpDsoy4Mae87n+UBFwnhj/TD
N8x6RXXhqZ69QC/AnkziN8DOece3rPb7U+X1wClcJKikJoY8+4IGozWuyF/8OjuLC785HLjiZWFW
52Mol+r83Wmdi29mR77dNJP59S948/wv03VrP4jJmaI9rTdAY81/uWOc2uNXVf9ya9T+R0EQmkdi
5m8Q1Re6QlDKjH2g4yeJoWcPt6AIrH3FUi0YFfiX+OSwyfPmmtSXmPd+2yFIRVo1u1QRR9EJBuUa
2z/H6YR7KDb6gpJ5QL9oW2K5QFOlDlLRGBFVw/rmqf5dm29cXz11BhRdaGauM32T+jgizyK2cV9B
wZ3dL+3xeMMo5nwZ+8wAF42Fq8Rz4O30Kx9+/UOqSwGWFKbq9uRM0Q7/CaxMqVWmUPD86sc+RfIc
rS72YkOSXq3Nz/+Jy9a1wFf1lkHl9t7EodwlyFja3I34uBufB1HNYLe7wFrLkpA7XRlLtxVAvhJI
7UAwRckAKiJO/wswyZmbzT1qmljSlQWMEoOhTdWKgWkB1rxJIKRXy5FBfc34Qmlu4qkin/GP0BI+
H7V7SNg8gp4YzCoSTaw+IUTfG/qP/6P5KkjClReWhNRJFyW6IVugMHQIizL0ey0pwGfIdlIar0gF
ov9b4xkwaO9RTmVJt9Bn2QTTyWMmbM8bhZpAek4mJgubCKKPsRqXNVdvFbx6N2gHMf4SR+jm9FEm
iUH6cYwK2KLuvKfm8rKqwPqiF1SGvsWtMNpBGILEi3TFRRNYJ2xu8sL6MrTrag2fMutqBZNhQ71H
bVXQ3GH2GqRl7evu2ebe7AYy0NPolzEAr5wjfW+zlyHIID6BCRgHW4mtugc0jf0eELteHu4MoVix
vx8S/ugUb0GspGjInKIeEIoiK5ISgSJOIE0TFZbJDb6mPeitbSVHX1Szrz+mA9UhuBdO6S0vWf/k
hZHpuPv9DMp+xvmS0HSgtvRf2CBV8br08gDBelnhQsHW3CzoFWrnkNLmie6dY+bAQX/M7f4niNSw
rzptbQ9SDJQ5eINq38uvW/PigZfRU+5HS6P166J9NTn7mwBD+U2s1ECsSoYsHjJtrP8uRl4xLEzY
GdWQb9GrBxqlVCnvbMd1F37hqLUHTKLsX7CQeGHiMVQP4AasI3UZVuQ+9ayOMoElqdKJoqi7K55n
WhGJM0E1Jgk1+5iRqPb+KDcf7PtkFas2Vx9sJXjF8FUeBJ4Y05nmMo8AEAHluIS4WdXFUce+P3OD
99GkmgpleDaf9TY7AlntUN5nu+1HCAjL2OXwm14CGySsnRZwCzU90mCfLFKjEOnoeV+FZ00c6uf/
4Z5nBBg8agb4bwVpvDblKhsQrhIuGpUMzhpKA1pXkAfSX+RG63HMZ66KVt466hfYTgjKDEpgMOKq
F8ndlgwsOtf+YJuV8VBvOxd9tOhptFLzwa9UfDkYc8S1BaKD+xb4JhmlPlM0iMnPKIDBSQwGy4yy
ZTO/+AtxDkWKN4N2G43fC4fMki8f6ttaeLUqVpqJ5g0ZfwhRDJRwHKxICJNf0rwPhW+u4Xtz8hV8
6bOjlroIoqTcCuzHuJUDUeM6TdDBzK36HeTt2DJcMF2mAxXEkPyJHCV/ZKZJVEVOwgWsa2kQpyXv
4RBGtsum2XjvAZafnvC01PE7eJ3krW6CbDm3AmKWJxQPnjA01mURk1FByqgxW6zeMHc114eZ8zMi
9bVDxXhFIs6M4SWGuibh64glh6jlyTIGoetoqbs05CySeieKgHYruAuCt0W5VNZuzBPGWes0l0D/
dCEsGRCpdRVSLvu01birXrM+iUOun+iTAwZBbZczTZD4wrRP/lPLKDHVwbfMPZWnXyFW/pVynPKt
QZe+Ba+55/eP1XdMqz1/iO0dry/oAa33UrOC9Pqtqv+MYif6fqMKhqHTqYPcVWbgjMthy3gekrxR
Am7i7j0ikj/a5X0yaqPnWfzFTQTsuqazPCl9vBDBGXZsNodv8LpQiCPJtD8ZK9U0653DyZW0COOq
OiYjWhHtUUbknzTLkuUPafQ0TCYcKDD5hNAMnWa1jst63zenIupib7UzQj5nrAC98ZXaJWN/AHQI
Jz87IpKk3V7fhbhwAdHviu858VkQyisUIFlzS6h5PYhxZm3WmYXtu0ph27XtuJok5NVjBRxSxjXH
V3Ci9oPJP7/EZnmwY+fBeBR+Ra74mbdL6c+MBxLb/bYj9TBNzfo1rdsBS0amVr8nNGp1iKlamjiB
8WNnkeEAPCcisF0+Yl6AhhYcvtyLPgdWQMSRQckNkymGc72OwxTqfkRbnzhxVfueyybAd0qlQhYI
RFKbu1KkpeMglNdOTDgLJz0uPVxyeQLTFu0/WhkGoczq7xIcteKlED9A4qa/rdoIzXmXgTWivONh
iybkPURUAbgrZ9idLBsIUB49Q4Pc+BCj7DsSth80yjGISYLqSe6oHVhBvOGEfZUCUFOTvzAWgx0i
c7VS6s5Bwa8mtLuDHsDue5R5T45tMDKWPWE2z0WkmyIMQirFOk9AF0pPGisaDl8SMasjGiJb9vbd
Ddq89ErMjS+j+2j9xoAdFL2lvUKY4N+CWXAnOqZY7hOKuqRv4mBJvZHW4KGrgmFg3VsSkyGiYiLU
TySVd68ynIfNVfCpHuKJZnoCRm8HEQ7m4Nr0mlzeM3ZKPXcZSv+0LdkbghiRm6EGOrJAH4/2peVm
Wtzvq0eBdg3T54aaxI5lSbtbkWi7nUFiDNYrAWEscIsZ8XBKH5hdhbKfiuxlFImNjJ83lrJKh4AV
GB2PaldixyCq/3qpB3jiMiEdLR5Q/gh39fVL3NOw8cL+VFtt/04NBegjxbAb2wtPDXFTx1pwsShT
SGOZTwjTRgiN39Mn5Y75DuhraoZN/vbxeGZrlOXyNgGd9SfISgIP1VSOeHW9pHXfhV4yht1v0lZ6
SyrvFJG357/HZZ41KX6ysf4DthpTb4ZT0/x6ocr09uT4/1tXmAYzSvx3t90LqiimJMYVWxGT/nnF
+88vwfIK/mVNFKaEoVRibslS7VaaCeqPP2Owtvv6r7zeuUx7i5gyLiIAGdnINofpTj8R4wpFaG2V
rRuNB9Mf7iyj2aRoFwYvlZkmR20rsbTiavwWMkOdFiX9LWaTjqbm58m64/xlm2tokElL6IVU+RUe
NZi0F0JEXcmJbe0+LCdSijHQnSzirUvuAEMAuX1c41Wm6nLo2dno5Af1wm9H16Lv5+dF/WOw+/rs
QAz9Uhrzz/cAibywW0UL19tT4KLiSgDO699HRvHG7w9h7Lhlw5FurdoKyj4gVOdAgHyffuaHWncd
TUurpt8ytRzJ6xLCDMI1Quiywkid3EPX9N/uWljeHJV0MMqNwRxfK8TAdpCqaD2x7YB5LdEINyOT
59fPuRWIEkUI47IHheFDL9+Y+EwujdRyfv3+eQUvAhd5Aa9273mEtwqZ/gSxlcAdZdp8yHXPhzAF
HBSXccsYeebsEKIuhvjYW3VA9mjyTrbFS03zaZnG208gtAA/N2+RsPGvsUubXxzSiS8JDQUL7nMW
uaM8dNifoveToeGRQG2kEIQDkZUIMebKcw36WcinGk6sd2AjdsyoOZDiXL1oYMdZH5+wb6bbbWc2
g1OjmWViCipRuoNCTe8/kdw2gYX6AnHWowCq6InqePQr7ZbebBXmL2D0E1hlUL2Xz7xcbi9ZiXwc
zL6GLVf97c5rTFcRnMatOP3La7MYYYfLI8oQ6SE7J3JZY2mIX/BViesLTbXFfavH1PYOflHjvFcb
NJGT6QPWa3QSv5eW+TzDH4Os6TQOYnbURWtIayqwWhZCDrqucSaEUP+uVlViDYLYP3uuVscCzRMy
ozziJhU45pPrB1sADG23+GgfSulMn/Z5OxQOIcmcoNAMTVObH1IqZzPza1RGSHMORl9a1Coc91fy
l9vbVMGorWAY5P0J72Amb5D6uNuN+r99EphrwtElsulZT7abLme227FX5jyHnPMUMkg83snFLtIu
/l+xv0Bh+WEaST4K95YPNC6d7llohBk7gcSGPDlmEuHUn9SPjNQCD7cGw4eO2WeTwX8KyzfZeji0
cpl8JIKbVsnIR7TOamMnnUWdrZfVnz960QRVaqlO9FVwnC3C5MoAlg/2p+4H098YjacqOLI4DZJG
b+CgzO4txkf+SLvgE+8YQEbHYR/yF/SVwz/wkBDJ1B9+kR4W6KcQcV3c6hnuEqIF+BVytetreE9S
uYUVQ6UzSmR8/wgNZ5zK0AhxmcRsEBtZqXlG1hjJJSIVxGYbyegMZElXNfxLCXw2Q9T1ox6/3vtn
AHbGTXPiYZM/nnD7xSvCzDx/oigbAqZktEshcjvGUgJ9qZOO1wPlilxOTCfdQ5xVek2vWvXf1lqa
SW8nlVRB2MyGLgYwLlwQxMVmN99w4yu44P83f9eux/moHVA4lOPMKJa4LXe13OMqZoB9y7fsDS7+
oZYnEtmhnf9t5OqA3oqCtHs25FbGmhjg2m+nYSm0Py7h5/Xltb0gPxTrpdTFZM/mls51zn1xCHKN
zr+Uyq2/lHWCsNxBHRHLzoam9eNuAbbmRLrCE1fZ/1onwvuiYMYVIY7s5aDlGAusnjoZ9uaLnjb8
SyjgO++xG5pZ4KGBGOWQWjGwjhkOofWFvJMYBwLC3u7ikFfwIyBIsdFbtbHCUgBfUKupw16bzyyU
xHLHVMs/SZ617fmgUQ9SLaZ4AdZeGJ2xnmmSHSdZ/IrvZbvHFv8TusKWDT7lxLdCQ7kuqnk8JMPb
5E1muvuXif8xAW8N6bBirX8l3wX2qeHG7nmfmbRFPnaPFWRsMDkG2Nz0LT16+vIxOWmUL/SSTYlq
HQTWmmXdzZUx0eJsS60dMbqBJT45qhYruMAU3MqjVabsrxJ3fwPHGCR3MWbaAFVlONPCjzEfeJ35
kPKnMWiRJKu0A1aRFW4OneDmBxjiXMPmc22JSSqQFcg0TtE5tC64/XiBHkhMYXMOChGJDLfJcl+T
zg1M5XcOxM0IdYQbwy0v7ywoHfZr9BtPShWMJn1da2ciSm4RKrhBcKLD90Ni1Jh86PhEh8u3QtrZ
1pmjLcKY1ayaYP+Z8m7xUqk3xZvxNcHoR2obSXrIZfjwAgs51gNS4IMzbt005thPtogN8dpHt5U9
kLt8Ctcftr//706xuCg6hLwG6W7cQL2r0NA6LFbhO7eGya7kWZ4zpc8rtRYnxgDS+oozUQV7dNS7
KRhnlAKL9s66hSu4FrQZ2slhu5eoYopSSk1bJXNblVaEH/nYjikBWBJKrTbs9j1TmeU0q4R8BAKR
/9GUcKVoFpsZW9JrLrw62ydqdsP10D/LFNYqi8ZfD8ijS2T5u7nu/KFR8fDD71/afZXh1/URP1mm
iN6vRmKmJYQH5rZizCdPFKyQlvWAbvPSaDSz3xHvRd0QXURUduLUHEnrXXp1Lm2WIKagX81lr/rl
cafRF0VH5xz4/oEw49NNLzyEjTHwNHCEqvJfH5+VgPAACCEOnyHUAvfCc40ux2rbpTHTnyt4c6Fw
xyHJSI4SZYUD83KtDHyTCZHSoZ1RTmjYUT37rUi09lOsG2apN2BnloRlUnu9qcdZ+uCXyb8zs7C5
bxReXUIhyYdSKIfol5cJYRrpy5+XoYIIRq+wzhqs2vtHeUp97XqHPkF9Z1HiDalHuqpx1EzXb7mP
M5xN+bRXzmm99Uetim/3gzrDUEJ5yPZNLB9/E2xoVAs8dr6Bxo1NKpZCfAgTjhIcpc+47GXPujKU
sJCp2BhGl9xywu3H4DgFFGIkkrgwiNj1JS2WKhXpzIspmCHf26QYBTMeBd3qUNttyJeoTOIvG41i
tw27gptIZU2ihywfEyP8dlFpvLMrBD9glUCeHRDp6dkgFePRs0QurL+ZaHTSqnWKtne6Ly4DKB+V
g7KxrNJcJJWT3JlaPrPckOfQz7vu4cr7PylPPZVHKopR3LOg/MMjZ5p8svr6mXQkig+u+q5GT52V
UP6CS246JeXVbwfWkZcHzQDRNNZqk+UFyzWCXrskJczE0xcZEZeNTeVuh1/QQ4MCmFsJ2n1XsJLK
oFxKk09LytQz6AKWiqbMH5QJqqz+TVRJrZP63h1LbF9euF01QCbfLCQjHGZCfAbfO+IugyTloDrY
D93qyrrqUw+qS40j2RUEBs1+R8JxELP+c//rMPqhHXuPaCjWA89XicPVLdZ/W8S/4Dctq/w+3vJd
4e3GhKIqj66TgH1+ZuJuHKltL/zpVpZwQi3WELmu91wooqbpf1Z5ekK0vnj6LiBYd7ek7FL46QyR
P3Kips8rvt3B1vMLmFEUx+LJKi4uC0VRMdaO0sZuLfSDnnFitpFpt4J1YBrgKo70rxNcxuXriNVh
YD4TiNXu79w4B19qrmVeH6dg6xpDTZP+t9nYT32bRLKtAAA3+Q6lsaCAYfEwTG+OXpv1H0Joy02P
i7iSJbo+GKLmVg2KXiTglhjYARIOnR0G4Eypl+17BUOmb+ngmoZpGKOZk0yospeKTGGFo9thIvLD
rtR5EK/8CDnZIblSU5PaBemqOZjwdnXZnxFTeosTwdHgN1qRaRFiml0a66/wOZd+KUo9g27Mbm2T
csOo6FFr7EY5r+8qpVPdEPW7aNnXWVVn5H7w+EmNvEns+7S/3YPpU2NwbDCLJyFD+nAVjAtbMoFi
eZzkE6JZ8x8q62oG/1eq6K0aEgC+cYZoFjEus4r1Vz36TKADO8HFWp1JKy8h9nn6Yft37mxLm1Zl
vnfuOZp2fo6YR7CDTYqzsoPp8U1WRE4bI5hX/dh0k28Jb9Mok3PpS4ABuH+8Nhhq0rRNrN0XvUU+
hE/vT0werqAU/M7qEwGASkTibJ650b3ovxZ94TbpJx/80SdljVPqVnw8Ge7e0r+n9m708FzKpb/1
4OrICZI0YXn2+OQ+gkdZpM+QL0y+LYTWVjtkMKoubTzmtrkafPb/G4XAYncrb9Z0aj3DKJOigXyh
z8mBjwGtUPoQ9gHZ5KMvPx8v3pbhJVsFM5zpNLMDNYJaVwhQIQftnDc5do+POgmr020XO2H9I3xz
UyIIWSZzoCU9aiqFGmlDJIbHtMvDO4dSv3ch2tWw8nfsSRTZx2RsoNNE75CwVsOB9UTWaQxJkMxs
e37rKbqLsnNfl5n0H/PJvq14/FSj9mKn+825tUfqI/Te2SQ9TtOugLJclNYkO5y1A9Dy2d6EG9s2
3isZxiSAsPHI4x+OMbiAt1nl0p+isq99NJEEoT0idtVqk6BSg1u4SkuDt8V425ewhI3tDxk3R+2U
Sv6iYwdQF8BJq6GQw/eo/kuwRvkV++veA7n39JEYN4qCe/Jr7tSP/fCMmr6SQIec2nPeZw7PFrNo
FtW1pc36uQTC4JyqnNHIm679zRAs0CpadjxO+0IPagPkM52i8j8TmovPa2KBucxr4WevfF4RvpHT
+vtymUQoNGa0/PE2V2S1qn2DzAqPFQ4xK1BpOS4tkVw39qA5TC+EYE/+Z6Ty95cUDmgjkpZ0J0Ax
RZUhDF/wx9UHzytra5YkPLu0REee1ednJaqww5j636zyw8nUf2VY7ajtUVVgHwFY+zcCM2Q5gtdl
zYKvZTlpjmfTzU8V+gXylD/K1aejnA9yliVkMjDO/8LRuEG/IwuQVPH3irkHIZ4lfKBtiV0JBko6
GXiGlRMcRdIfplbTKVwLJaV1tGl4SHC/UpLdUaE+unt0Fbu6y5HwFYCvd6SoJgwChtaQQTgVM//p
4GAIq+gsHyy8dF7lTS0MsnjPiBa7xHHD8O7PCY7qbgpCxlSqGbxdibvejVM1E6DRQ4sMPaaU0yRl
lcVhEcqpRVLisKSvMBawflRl+ZjiOgVseG4DAQY3OYkAina+n+nJ/MGbQMhqY/+NYxkiv+XOQygZ
9BMQwkDJvL45pe95WLE3+HpTv4L8ONhb1tDY47jlbayA4+SlmAaUcnRz+Jh8Hf80DbNLBsbBSLZz
mwtZpRj9rXdfZRzvcU13tJbmvNMZFRed/Qm/Sfd75rDiX5lEWHNvR2s+uFPl0b8LrmxsoJGpwxzu
eMDp2Jzq/ac6lNNxFryCtdCFE1llTEaCy2rS5o+r2p5boEB22Ik5kOcDE/6yhfm/FexNHzrXGbec
L8MZ1kRiG5qXO6HZKTOifuH4n8Slx7g/BbF2LmBBwpSbDKj6TvzQHiK4ta9+OZOym8OdQX40yLpR
lZK98mlc0KbX8v2ONxp3kNDbfCyygyy0U5d3wMJGLWfevoOcoxcv6DI0b10yDXLI4/spU3bUi2vv
GDSq+SgiZYscx5m1hDwcoyzn+aNHdjzh20E+9GOg1GyG6KyXCXaIjiZdS10rq3cRebTT1coMU70d
BRjiGyu20rbdnf2zuUVl/HuHKRn+tFDMIwOboBFBHGIcClyvZM1Le145RlGyfA0v1fxop6/Z1jSY
E8CtNXbN1B6OZN/t5S/dke0exsOew6pyfWJlPCVo3lA1bAHJAM8Q9bVMS8XU4bJqdy7YrQg44Twd
CY79ilDbAC5q/Nj3KHiGQd+TS8EzDTmDD9nwmm4GEaK9EexhCR+XYi9cBJbsn9KiP0RgQbFjY7wg
7cBLkgjZkNX3m5AJQUfpr3qegiro0A3G09fce487tezS8YJ89mI6K/r5VVgFh5jvxxXBEvsZgWSx
R5HGPWPF7AxQI2CTsSE9hqUz7yyEOvLcEj7yVZ9ul1tjDN1qh2hkLKMwtrR4T5iIFvgFquJAEChD
K5JJ/PbUqaG6kXwyHt/5ldp1fXzCPU0H71jZlI6zsHIwcDoLSy7wikoJmMal9ybFsJyCZYh78UJ0
in+Dz5lHlZor+1dEQm6uFVanfhJV7ZjXIcqsLbqAmfgAIrxhu8bAmetGuQ0tSDLHoNJ5oFDX1XlT
gbZ8LPye64PtLxgFriWZCP/5+sXrI4jcuQlf/WkEDAAOkcc7aYF8x9lUI239DCSKk3SmP8IZmdZD
pSM0Q9/ChdT+eFGBUHyV9dnuWWTQjIk/kJ9CBqT5M7Sdi82vIMmpQ0IwPN8wGvVg2MMCFXPHpZL/
veOR2smTy2sBe646i2SN4N40FlIjNj9018xLWGSOkcsG5ueHYplxvixJykSJiCB3TqarM3E0wnE9
9PcTUj82GOUGvsGazzHL7vnzEubl3JGZqBFqYi949S8BmA62rGCkcCXm4hNzlyv8GJmSNXhUGC8B
KT9VTlYI5QKm9K4r0FFCxmwnH2tEO2tD2Btep+st32U+S3Tu4ZLxZIEDsenETfMq+jKoZdYO6f/4
yY1GtOK8iL8dMrnmalKUkG8JLecKZutB/xBikB26qqobWRQ0B6knbT+16caqdAERd+XxauXHDX7T
UBJan2WJT7iRQQKZcpSRLh51pOosxQEyBvBdpoJKmcLb1Ihom2+TSEx+UBZORl0QDtuuM+zcKGqM
WwjtV56eprcKJ7qHNv1Ex+1HkMnF+fMWyB+i1W9oYu9pIHCYgCcOFpq9bY+mi/JgS1p7ad55gjvg
UgXGttYy2CLpOrzlVSauwl5nkSUiH/QP7DZyg1lciHrqPYH76otAH4fS6hRs0Rrzc87WG3mRzcMk
xgY7hpLgakhYJuZzL42dDPCtm37g/SnJFP1LxbgYiUJK6PPNAOtmFmDsjYyHZaMROvEegkirphuA
GNWayjzT/+aecfI8XLn+Q4+o8E+gnFDQDyd3qenTJ7Joi0ZSprAtG++FQgg0P2aIyRTu59uySIbM
AsIW18zY3G3QuNcRwU/QFWqXEwKHt+2QBCfQa6pLMLOrkzMWrzSPrFqGdsRtJyojQ1vdMt7ZdO6t
wB6nHtvPCUDNZPeP3HdZQ5YVayNw6OFOxPWU+jbGb+kro79bBD4/OGsRwfnDzPFdMerKqGE60fHk
Om4mPyQ6XjDPQV+qw+dpfacKm6Gq/8ZwgKjx2D8MnWEl7jdIDYcxtoxmSjWegvzs/HXp3pawBRAm
yGVEmtXlIFImY8FX3UBY16/asjX3P6IVcgYEHShjJml0u2tkosMFMH8vdju0VBqJxe57YP3sgNbr
wO5u9NeWsSyVTCx7Bmo1Om6JRET7m4J9zE8+1zygxqdqRB4iGkeCGeW3g1sN1RzBi2B9Wc9qnw8n
WPBebT5YuQNEd4w1E+NKBscnVRDkriQNTijpRoRqfjX7kpsi0knSXrDjLUJDNEPBbgZevyHE8CXX
Fnjx3CgIZk8I2rOtWiBerk2xvg+Qjan7Q8e86BDYZP6s+EIxGD3RulzEiLvx/4h+plhUxVo+lOUg
5SKSPj1aklz2ZAZ0KqQzoNDt+W2cWGVvjdHNWsQiLqBsHGwNYYRWjdA9ti/j3C0qp6MHWxbyjzqj
RO78oN6T3Q2QuhSAeyRdJjxwjLLYLL5HSCxUf8R96mO5NotnLt0V7qWwtd8bAJkskNRe1GaDLza4
Dm9PK+ea02Qe7wG5Ci0Nt3xL2UR1oZzP4WXmRaNFmwjH2+gci4sIypbSJB5WA1m7fasLDRpzFezX
bhv96yG42g7fQV1T/2I47ejeDtj/FsZh0JXr3X2aKvzgvkUfRJlVTDTxA1H4o2p41CrOV9uuKfG7
8e0fL/XbpSCwm2Q/Z/iVGs1V4xPQtNfkjJYLv0NkEB/uFn/7/pqFmOAt4l7ErVaFvmmjiIMeQeF0
wxVwvL/BXjTCbBerFEZC4cynGmbt1FzvNY9MIgn6gNosA1OqBgsuROTERP4nEYkn75EsXMoFpPEH
X/wPA1tQ5640tYwbg9dVKLzaEGTCSw1IBNe1TCxhOhv+LnUOVcCECVN0oEcRDRuyuuu+8OeiUGMN
tr8XxVdzMF4HLy+TcoqjwzZpZIExV7aHbGkHQU2BcaasOx9Fbv7NuP/dv7H7mSH5jvSJgSQ0BIYf
hFN8t35hqo8ltVvJMIafPjMeSU6zZAa0jSk7jArOG7LjC+I/X/eo7+pEA92F9pwwGbG93mKe7ZJd
IGUJCzTjfDwIxO1ja+JatYLlulutOTbmF1fj9yGB1zTQlJR9WONZ51o7Y3Zk04bEkK6c16XasjxA
FppGEtjK1HukxKAVct9AUYMy/SI4/nQzAMRRJmAIfSsiZWSSu768C7zAkkPeo3j+O6zVmKazy9yt
3jHAI87zb3IK1b05Qm7VPn37CGX/fY2y8k6kFBU/lx37sRm/IAIhup7B5lBpyIlO8ngHGbz6WFao
1uID5a4P/iL0ycpCMUCb2zsxIth4RMjpZ8kaVm2ZqBiFrrxBbj09BzjFnaoKWb7qXAD8I0E76Oqy
p2zKU8FawLgxqExQ4+jEIsHacZqXZ69IHaBYIwWBDZM2KySTN1aNImuETHQeAxk/az5KmXizrcFd
Sact/e+RRQgpMlb9auLe/RmXn/3StM88gVIqYQ/v+W9zbD2aWx0s2kciASFmrkKCFfUp5Eorr2ix
z3IKSt/w2fTxK7A0IWYg0+Z0OtOqZy9UG8ymrNiH4wQhNclDD071QG34F1GyB1dvm8LvwUcCdEwy
eEAXfVSdKFguBEwNNyIHHPDUuqVFvep20zkLEatozfdz/xHAbZLP00fbqfdc78tXjaW0LshsMq2O
4BJ6G3v2XdjzAk54ph07glqDzMGAnyBfx3GVGiQRnyH4B+2lHiA9HN4yVgU8mDvie64+XM2mM2gj
D6KVwSW5lvK117d4FO89ZQ/D2f25m5ek6K+xQd/mD7ELEyeLSJQLmnuvQzfnXI5D8w4vW+M+i8aC
AuNpuIoicr9R4dMD2P1kJwcYO+9rIy5BbHNKGd2R8bY1sct8BHNl/V0G8sLLMYXEr3WIJeWM8ev7
xOoTwAfw2sEv86zuEEOatKItt3c1DEUsCeUC2OfNRHjX36spiDiWkm+r5bqMlm0VuCeVFmFqCDH/
lZqiPBvDpupzZAeOCPvPoY9iDycFnKbjef+SLfummZ2GXXdLB8ecf3WnW1N06FBar/fKQtpWXacB
O1IMCuq0JSmPbZ1g/gMP9cztQ6nWLJRAb2T3IKc5niYT9XNmVO7zxoeibbQuYzOw+Hdd6bXXrcm7
xZbQ2NbGGFSNFXMEGImedNtca9THIL4FoNdi7jGuenlQ4dxvX/a0yRZ+k4hZAx0XNrG+fd+RsmiC
mdnQ5lxj5jJe4qtmkJ7R8Wx/a8r5jn62OFkKUNTctcQf/4Km4GL3e+YzkXKdXrXn3B3gcaIvNsuB
bsBg/4K1clfToMHEeGbiATJ/kfG/RhIdOkLy2c+udBJfZO2AeWVKB7I3LAdxZ5K24pJ5aekcBbq4
UiinDHe5TL5wWcdMzSvQ3Ur0iOjSmfv46UE2OB2ICkWyV46j6+PnnkXpn9tkxgH/fsaXZsKiiwjV
5LxwgUSX3UM9cC5qPWBCIgl15NHCh70ar3XCI2CFFtU0x8Gp+BriSKk7Ojjng5qqhTT59l06wiEX
8LbGv4dnfFJ1KS+ywITC/hvEItkz9R7X1psrw2KUOptdP9JHTGdDyC6ijApWHRuA7gQF7NOAwuGZ
GZ+8gXQKEDeXIP6hoBdtnMGJGS7ApGXaddeybnmCgIQoPuZYEjjMyNs/XulzGri0Ohx7iYStIlwZ
Q2k/1B0NS0l32FhZghNsZXRca8J9rcEYQLeVd++RYVnjFOdla17634+riBIywUQlNseePqK2QGkf
O5ndlfJyPdv9W/zgkdHsTQfXowNP0Aj92QLv1SCDCIux/GU0urGVVvKwI+Si6qaYXOhIn0TE7d6u
rhMZXWwR7ILVseAaRZ4nsLmA1m/FIOzVJ1cvfbY4I4g2OQJ0cls4SVXfzt5sqYAxpia04DDhC6mT
C+46A5uDn48l86g18i1AT18LktvTSL7+aHbuxKTMxVMDrNYPazbzSCuqSTAY6L/izR8sXfhDvBd3
yCwNLS42vDpgPvC4j26SV+atUCDr3yCdK8YVnl9XelGp0/F998csplEoStDMg7GTKQHLzsYsQUnC
hpAxsESReOEUjbqcZvJDV29Ih1G3C/QWeGea2m3K9TF9dcnVIN8iL+ZBIEJ9fMnG3uPPZ+u8AIRR
UG7ObH7OFn03eVA5KhsXV2qefjzxVNQZXTz654rIQMED84FxW1ZtLRCh4Hrk4JCPf0p/dTzqxYtn
v84VJ1CGvahcYEIn1GvxEOzVWin80280DO4rzpuzYr2ZSdgzv4Wo/W2ApLZ/gi2Ofs9KOsiv3v9Z
GB0Pxf9AeoGLNh2lnxdvRDSfQ4kk6I2p+RI/2tKYwvY9nWsGWDX6Mz9Z71Hn6tH+Vc5TMBpQ+I8E
wZay0rJ+2lLV8SmRz5uGrgwBh2GDEndeebN1v8w0HW02CUZMhUZn8S/O4JDTLLOgaxbFtp+qQMta
8NU5SMtWNnmU6y0Og7qIMAulvkipZVV3AUqL7lys/iCXHsuJSyBkb2KRI6GSKvtALku/LxJIJ74U
M3g+7kUv6iP1HYTsaSkwht3V5eh6uoIGB8jUkHabQccksVDDOi7RgKFtwPoM4QN85jlypE+5JmyG
VlNQlC7LXsSpJmiFl0qmkSKeZNFKaIwKJyd4NjJx5vAYjC6aP6OiI9RHmxCg9Q7mQJOG6dhYc0mT
yinj5KBsAQnQ3oM8mWRQqPw0Joseu80NNRk8zkoYvEnF8zHI0gpf14fHb9ZZ81w/vQTUv/Dq0NnN
nmPBM7auTKrG+h6XzGsfNKgqyk+jGdnWXq5vs3p0F85cubFRA76GNdayFTfczG4eF6+KRZZqwaln
9JkGRY+dIjsZMBLdth9zLjad9Le01NjDYny8Lm3vR2ioWSqRdzCJhWEQAvCDssks6ehcNUHeOf2M
8kBbt4jcsgPKNA6OHe3g4NhWEnu+ezvY9W8osomhXH78luf+9OsTYavHx/ushDwsAef+pBz7RkQG
hSRa3COAm5JEeRgFEXt1EqRse2sQaQCOXQOwdkgIE8lnwW9DGEInWKl+SCy1ffnaPhjqJyl20EL8
C0VNBdYt/VpnKRMc2ImRmZvdzSGR1ZlhZwwBM+qtvgHO3oZVY1T6ifMnol13RABzqMJTJNnmknON
R/Dd1IgtpKC+Ux1D5dBcNygs0qUXeZL6AdewRG5ksHzVJQlBQSrOtO6GRPlgRqveM7gCMBOIBPwp
C39KvvT49hxxOrzP51Xpokw/RtmqI7Lbj5AZ94GyMSn+TYHBp/nexpBSBGfPOlj3BAchIYQ78pVv
IgOwHjv5XewMoE1iV1+x/AEZAoIlNu2LCSdnTITesqdgqPYYnuZGBE7mVdnOcV3IuvKcHo/aTAFN
niv/U9xV6OP6aG4z2gaAbs+OepChGqC9Y9FnepCVJZmVkWcDViE+k2LohcbIfMnYGZNt4CMS6OgH
CkgDBAK37lC+Fiq7uJ1XEIPFE9bXGQBk2DHQrgDmivrjr5fi0FfhHfG1PKvUkr/ZCqm8VhR56yqx
wHEd+uRYslx9mK/PO1wi1zRhITsRPt3iOSZXMEsKi1A40MSF8CFhfv1vlHFWeuPTlK9v5GM1/Tjg
lSdvlY/Dy9Dc0AsIFaCL8AzfAZ0xnDdunLybXPEncUZRpLeqoGekTKHXZOWGrRm6UlPIFE0BEzBd
+c62D5Bo9Y8WMYLOFumjV6QIq8LohjQcYyUdzHwvYZ9j0Xw8AF+dUDtOs8I8eT7pOOJJ+12U899w
Ju+xyFNN8OYEGLgKRcGbMQh9HVo5qijNtOO8MHL13YxlvyS+eDUVmPVy584f3uTTLFZdqo83Y+zt
2vmn03gXTRix387cVVUzxruoVFSQNDGITEk8CN8gAYvAHEQyrSZ2qjD3qJwmQVoLwIUzZYio2+Fb
Gk+MyVVgSt/K+XSo0w5l4pdNdb3srRgFjt+BUuL4lqB5+R6koCf9rAA5YqwxMyayqdy2Raw31I+I
StvTgcZJ6qXEsK3H+yK1UZf2YB75c8v89n0BJcTOxx3rjEyU041HwtXkXJ1KzG88rZY5qpd+bYO/
bkcx8b9j9Wx51tHO39Py1h+Ry+1YnL59UYae5BdOAbrH4qFn1MH6Skq4GlN74W0xhpf8r0rJymCn
cgUBJyHX8w1F7LKqCquaDnZ98iBhRyorNBPE8tiETc+o8/AauQWSpi/aNAVjTJKMxZZF1tb+g/bd
rW95DP/Un2xx9YaocM+SI2Yg6jU8NGEh2JPWvy91/XrviWzB++DbpNcWyd06Zgiq592BEsZz191T
mV0qL/WHK+mUA59CWJUcQESxnYKLcM967w21fNLHrGHORxo+biqUJLna7SFdd3azuO0fFvQxyF8B
ln7Ti4aU7gW2YhU6YldxbWaE4xzv2ZUNZymjOmYWDgHXoVCmSIBBPqDD7GvZ5dqVpdnXCa2jBnno
ekt07fFyo2UlwPgu369FCKZKxZEK0dHtQVNNFRnRzDK6kBwl+nZ0RcZbifj6n1QIEk7HSt8SAU2g
DSj3TEQuRdLPkAZEXLBuLUQAZguukCK2HoRvHKII6HRGDcDpw7zIjY2UKT/p/YusBxTxHtP/Uc+m
yWScJ1yVRQiJyOuGEUy6TljnA2bX1r0OXD4YN7y7cqmn8gXd/uSFjI6dDJZzQ8YX/O8C15Dd8rtK
LVWYdh5+lOc02H0lpt9D8mDGfKeLycx72UWdpTC1U4W2D9qUTu8dwyMTp1E7rPg5nj5Puq4jYgNM
hYO52IqDmBkydR2eKFITf68116qN3t848aF0fvVP5WWD6XwRqKcykfKBxKwIpD/rqGSvlU9dPGm3
Gbwf5pTQ9tUAx/Gn97kQ2qtLahVyOnWHaOETpm4Be55jiFCBDmD1BbrM7sTjCaTlYfsH02+akyOT
ZVbqTNnTBPuwvKcWc50TzbHuzxi8QSavcpuQ3ywLacZ/WbtRdM5Jqgdi1YZPZd2r7zCss0hLRvhp
foDx8yHefy62MlUes1sQT2w7H9IGZvJHtPFle+GeYpiQYFnmgTc6SywUVnUu0lGWTemMCPkER9gd
inVFFSKTUTE/2frD+AQPf8epISLjz9EjSghH8ou5wGkkBqy3PbramMhQOj//m7FDMSZ2BjZu87/o
N0MYmC3zI6uHYwlliM3+M0ZOHSRH+j5k6e5r26v7KgTB/amSsrke4y17jp7r7FbaEQVcTZLS4oat
p+v9a9lWblMig8JqtF2eO/2chV16YK0wQM6H4bsYzdHg4VJ7zWIufKJMNeFIUKZrAqnSQwOBz4Vi
cPPHDd9LnvvkBgiV/3UNIZYi6YlX4Ev3UVQ9fSHQcsPTDmOXZGDyTx21F1FMNlMTDsXyYmAgqbPq
rlOIderRAOXqrqg2VB7QBT2dXbQYMtK9+W73wRdvKEHbQFHP0qlcN0+9+hvx9WTgnY9O5mUBRiGC
PM2eWO+nax4sUxPnfj86mFKWKGOpEGLB9uLJ9V9gJCU1KBPYwoAl7BEUZCF1lfv1Hsz5JNKLGmVW
1dEwZzMlIqSYvYipSak0mGaiOFiKfFQh+DujOY/6FiINajC9Ns/OPTf/JEbLB3II2+9oLO/4dH+S
X76XZHPMc0N0YGEoiVGkOgRmRHyXvIDhxs9fWDJh9THOi9lCgv//pvJPpKxMSRs4lOyMO3scFV0i
HcV30mdthm3idrrJOT3t/RN9+BKHb+XBq/iBm7ig4RMBRhzK0yGVI2wcZkV5eQ0R+00CxEPfIhd1
1AsToEflpajTmfF/pjxciWWuLh+F/CMz3F/gGqobYKAqOeAg8bXG/osVK+m55hhysl1maiTFkfLT
Ol72fcNaoGAJ8nCJjCbDu57vfWKHJmqeJTksV/6bbqsX5eLna7suhpIWujuzPTgi4AYTF0Ick+7T
pcdtr083M//r6DCJoeMS0+5mjom7WoW+si4nip2+dst6xILrWrB1lSnau4LILYIJPgeePWDh8+b+
358h+b17OsCWDtxIqemK1NmZUqzlTX7U7BaP8yYrXzHaLn/zqnOMH99zNxDfynrUCkZ3V9vzq8t6
Q9LzUuW+lim4CyoeJ/xNwmf/bP4vRRaZnNyEnqyvlrIFMI3X2kl5n0Qx9n7Loig9g2a0F2Xce4UZ
eX3gR9YUJXjgv+xJA/am1vDSAmnuCSNL8HTTVY9CzflETWfyT9x4kglB/f1pUKP1vv4aNu8xfwyT
7ZKjONJoc3uSxafdJXE8BoW1vNOb/Hw+dtha9A+3iuDHCAxY5UgxYG1G1rTj8Dyu9nVUS3fL66uD
roh/0eTgxuTC8/BsVRRjUyLT395iTMFJo6fsHcBJgJjlIqNAAQcLhRczhNp49zKe2rIbgxZgQkVJ
BRxlYju13iHL2ltAlqPnpGGf0WV2o5DC6BzGzOmTA9wuR81UmqIk1tWN/kTVxc6sjwjIwD3yhv0D
jBG2GNDlS8CsTmx1OMrs0WH6B3z8X+MqDXnT3H1SNkKRSbCvJy+6xxmYnhnrDExtF+blGn0KEpuq
pRHBx3ukB1XvNuYEv4ryvrNDdRCV2WAtgorrV06dyRQdLUbEAKljSIkdR+UQqoQhGP2t0XMU4Wct
+LeTccceTlZx2ThGwyEDReKtIMAjNCKyUrCuYCx3xspcgLnmsbg+Efk9nRGYy7LDbQhz9LYoAwE1
rDDHdVgq2OmDc9H7uMRzVzwHciy9EcjJgV3zb1wiA20fQnHqlnQDRFhtPEjLFswmsgYruKul7baR
qt823y/hBhHGvNKaMKGu/c6zV38H69nr3MgmyJiH1N6HbitBRcGQCaO+4OCFV7fwl4qFF+1NNo3i
u0Maj4DoQvDnoJhXszmapl3ykYsxbvnh88hLzJiTY+U6mRPTEzmFXZRhdDECGY7pdn03Id9SXTwq
PiryOaTsrcnNc+kLgcbSCYHa+6Nj9sRpsPJEVjSLNywQBQMiYOROGPPvxlfpuF93NEpnprGvT++f
Zt+8csbPcNHULkbY+LBGuA6AO+JaJhkJoJE8Fm4QCqFooOxdcRVJgcJDhoGtxgZzxgBkAm0XSYem
sKXXHp8mGoYEDe1ZfjE49oGNhzWvZ1zgAOW7DzY7RXXZbj+biv/1htSkDfBFFkoEIkcDuKR66Kow
0rRQ3NzewuFhhGRpqTQmH5iD52Geq6dyk9Q3rPPsd+hFUfNPmCtcmqpfxPO4Cx9f2yyEwBiQzbpi
uwAprOQKIdFZqJaCWeNJm8/v+Uac5rsghls1bFlB//bRdUclzA/Bo7lsYM7NfwPDks9A3EHy3l4R
D+EvLAE7xYLfzSA3uQ0jJ3EK3EsWyp7nJ/m0Y7cOEh3QaHP2M3s++DTHM5hMmbPzyHnjItDKWQ5N
Op5+otEKjxxUBdmWhRlD7OQ7/UIbL5FUHLCBNC9yqECqqf7JE5W7rZbvPaoX/5BIAND1n5dYjWq/
Cm1XjKEZd9pxlvizquDVI9rlpfQtrUi0AhaSEL+/hCf2UwU4V15aa0rRQv54FQjn8Q/OPQ/l3eFT
1+4u3dByJTlcWd1Q2sIWMxF3Csp3amLfPfcJF5JN2np4+J/hybS04jvDh0TbwIL6Kee7PdCL0jMy
gkcmC+4W3d8YWDPj2sSUk6pJpH+VI9zCB7vDDeUQkYNLAceIQXIp0Ac5CdRYxzvLolgtx4JcLR0x
ZNJA+NtehHR7PTK+gbvm3j/7S1uLj1ra0GQIaIir8RqIn0SyG98qThgzg7G+doel5v8Y8hP/zsg3
+EwzhDusPS6tddhjEIvstP/rszPMLj4/yc7UaNsDhZt0QGCPAZAg4nUMF/H0zIpYIk6i/VOk05z2
nTGqbM1n10cHf6QR5svYhI7IxnYkqLXzdPkYW2hzqWIPl7mZQqX44nxlrv8LY8P0tOSsPpFV+MGg
/o78YwHgZzfQngSSsTYRcaJtTG2HdFW7R00kJ9XpATGItTpWO0uSO4UiPgkhIAXbxDxctvGLW3fX
kKJC105vjNdRI5SDi94dzxwHtk3zuKDby69XyWwvdVYTe+mxIl0Tx9vcZhQ/EI0ojfR20wuEubXP
LAt6r5mb6nlsnFxPwHmn0OvL7HuS21QnWQgfT2xDO0iJs9Gu3+kACR7XIIqxoiAv+7UYi2wJ6SbV
vwBtkSOPYll8zLqe2Q4HKt7JT76gaNnOGU9hN3yIaEI8khlr1Ft/jvulEQ+WAF6K/BDulz5vssVw
Ed8Xm21WQBIcXm1Hkd5qpgJbvZZZzUbVaeq8qqM0jzQZ2DDEYovDdIphOZvprUF46Tl//U5NGdRS
iCrEwnIQ8r/fut8ymQFRBxGSgdz0vlpyDAnKml3qs4kcz07B2mkHa8Skl7rimn4ALDiIvVBkd1k+
Ae4GMVaeGLzkdGXXpRdfaTCXAe18L+hnXsEr2YbCf0biNWOL93vJpSnVocVHJJbM5y2evQEGMGP2
gni/7jjlrGrN/LxVoA0Lxdr4UgRnG2eQ3fjbrM9aF+kXnoQMjIZtl22ld5tieTrvQ5tJyTl6d3Qk
6CwNr3fqe5pU6q9eGUbYZ4/EhrkqqzV4axRPfNQgY7Glmf9WVgC3jSfr1UJAiC/0iaudCp9kGabg
yc5QaNTe9ehv2eiZ+5e066Ho1BCXHFGUWC/M6SWCYT8hhK5yjN56heUx0YX93jDrykErZMxamsTO
54FK3st4hk+dXhWrxKgfjgKQPBocc5DIOV5ipAsikJHKvvPd/7RRhuJD3+iF13mgeBmSLvwWbTd7
DCBUWhigAxMzFSzv53CQh7/T7Df1MFX+W2w8VIoaT8yHooCaRRGGuZOtMb+cVEoHj+TyL0U04lep
WTdXTk7obGmSYQ+n8mSkkeOFmj2iM7NMMyKuxw9da3D89qeMOg5gA1/opVW9JvmPp6W+9Ds+K2Qy
FttKcDKpjhYmNYMFcjov158ggWsokwjO7ZZm4Q6du446yU4GJr1BGFyDUGLxgIoO9Mtxi0eQpHnn
b4EEu6w12li+3HgH9w2ivX6SaoUIxvJ+59B8KNkZJrcyzrMN/2Apq1kfs9YQ2BwE9TEz0crW6KQv
7GcS72Qnl/E6O9NYmK8c9LtfNUw76zg8Y32AOnrHoqGLqpao+GzG+QQShqCP4A0Rv/5uc3/FUsVY
qUlibVsc7deZIY146sxXlB24ZqELb9nLJsdfF57c2O+DC3ui+JUultb2sMbV7kz+XYRFRwUjLUfi
fqr+8a/0chY+iqlYv4I2nRjvUbiz+m5NVRz4SiRcQ/uzxhv65KsLWDALkXIRVYPw2UqTMVboYfPZ
827dOchD7O4V0WszoUdtxc7JFcESUqfHLHkRdJGkDHJjac3cGIp+xRmE60LKOgGVy73rMzzEsc4e
gGOsCLraB4GP0wLBvdRYs7ufqpz15NyQUi5b6CDuNhKcFyfJboJHTSOrBn380W26Dqv8FztfcWqn
xiapXaomXVaNeBcvGMu0sI1arz0SdNW6ZlSnJocEGOvnv16UgoONtTZPcmdVZzam4XNdUZ5NYv83
qo6wKdyGhjJ5R6xRGtn8wJhIqWzhF9u+nC/wavMNXFAoZ1tJFV4bPkeBOXIDOGIyrdBRKQyo8kaH
txDL638N/RzBUgKIHusDPfM8ho+HsrqZAtGL22gcMh/inoUmV/FYySTvkUWoWGv+ZwCCKIKBMH+x
kJ7yCN/GKu7PEN5IAXAX0rPdOzwosRItHTGJDCFHZDFqQpzgdLPikFVf23w00jIvT40qi2v68db3
WZ4iNAcjof0R4hg+3atWH97soo75BFmxeiWJJz+qsCu5l8BOZ1LlgTB43zxQEgg0QhxzYT+gx2Ds
rfYdH0iomnDG0hJVSWrEjp/+KYbHbWFb3whdSU7sR7BLoGv+mSWB6iA7H6bb1XRepqDc4uTBheVD
EFMQx6JvfBzHjSImLae0XNhvTriEprqmkRAeUzy/QhuJAkjdIucScmg8gyy3LjsWE1wxRBKWkUXM
XdMtntaRiwNU082sgT38QIxdhJOZ3NU0FRdz6mHRpHvTgUg8OFbIuri4L8GSCXKTsp5HMfQuHsqR
1ZouLS4rYR3Ap7a7oF5ytes+gPGFPKb40izUsZiUYGjMTbJmmtyZpwVpR2dHbxKeUTVZRPOpjcDg
CCS26UfduPw6Q12eax02u/CnfpeNrt2jx7I8MkbPfAU1lHxsgOwaPhSO2XAjyETQdynGUJ0rjM+L
kpK4HIx2vnMYDZjx1wX399aUDM5uWXse9WZ/k52jYZsUTdXbMJyQNT/avwmptOFgj1PeHBM0IcTl
bx9+W6FHVhUddC5VCxdjqb2uMujPFTU9KZ3ifqVpiC1zW/0Cmsung0dBXnpBrTNM1Dfuzr2fm+40
sRTXhdsbM/YbJJ+Qs5++c/J59od2rxGEQPPwmpM7RBZ8h6Ppe5gkQpxr6lA50BUGcqjrkOp/bWjD
Eqbw6eZWbD2/iiXQ+VOR8u8a19rFv98QvTS7OrbNs+Q3bfLO8xgqR0nVs/vKDv/ehYGzXzujg0CT
avDhLZzUwquxn2MZnzkrcfD1ADBOIVVRz1UCOjkJMe6af+rP8/wNmGm/MECjGlxn+SvDbjMJePCo
Vjpjb94kPk4nRjsjiZ4qzmkNjG/dCMHAvzz9A6Co+RRGOEMZRyDprXySFWVXe64P3h0NvxqDraM1
PA3CUVerAD/6ZSwFZUbb8V998/7ytnZ5QLYBf5APZJ26YNeo3Vxy9whA4Nmh7fxtpMzZygzIyTr6
BBesdKAoFxIsIrq0zp/jYbvFqurMk8LZ46qTd9Wr+cHVnpyrkWrFXrFcCwl3EMDWHbpGK38pG6B9
xQNk5NvmOHyxlq1SFJgXlhmDQ8xutt7wDFrOUgq/bmB4UMAHtMsSjfhTkHJIVNSPTELKEEHfoZ9B
tm9bcvAdpHqG0Chf9IQ2TM7t55JsSxB2QLIIWtqVbJq6VHhiwZj3QZHa6OAOwPbmTmpP+ThLuqQq
VIUgqnO9prNO1lZWDgnzOgB47lS0yHj+JFXlJqc4Acbo6ftzYk8Xr7Ccy8lten0QHIi3uZIUNZt+
KytQEwTzKP7QUFbUiVBtADJkprptToJMgpqKJrKvCpzFir/8xe+z08xrQsHmVKJWKRMaBxHxzjOs
Vs0hcYUH77fcsKLG01MS5XYHvLAOkx3UF2bHC7niSaRUFo+zxRdTVZPtgxbxCYVlyqw8hm5B8eP/
XTF28P+EM1oKrNVh7ipKE5o5bgx9PjvCuIpJnP4TCmSdpCH9ZBhBx3irbsP1Xq5nY1Vtnoa2KoFT
xhUeH5NZVN8sz+8VZa5CW2L7lxvQyMbUMjawnSbjz6YkYmmERBQbCJ9Y3MsS3++fA+OPDfvYyfP+
NN6lptp/yY8MnQ/h9YJCfX46SrKIN8t4E5gWO549CFOL6ZbFjj5UQFZ/L4tGA/1l0cGoyLOUQPjT
Stb+/jJp9VvB37CTYkN6xCJsVQIQKIWSixT5SDeztYbpwNNjnw4QPHkE0lAeb1Ibeu8BqEXH3iuF
teQXr5wWXcw5Okq3jfgy64fbkX5skirNiOvSXR164b3ari+LeKCQV3KTR4ABtd1sWls9fTe5cvmE
3opjiauGfoFATiw4ZFMPMuEVlhS8/Bg4fE+i3aOHWH2quH7CnjoOyIrX+WVPpGKvvBPkKx09bhu+
BW9C6AopPbdOytOzndIpm2g9t2OjmTteLxATqOSeGfHT4JgD6D/wLldNjfwzuTsu+wwjw8ewnLYJ
j6kduPGZqeDR8+f3jseW83k3mfp2P9yXzUKfS9kyksksiTR/vL8oAbLedQUUOhnLlCoroYA6ftWN
3ZhH3NBoieBtCjuXk0PXGv/ZfCc+lQwcPoQrBCbohWFOLwljcrFH7lwGUAYc090cU1uSimBNBW/e
FpYK3dJuyHnoCpnhhXQwOw7QrWkgzZYZt9+PCRmFxB9is+TrWnIgyG+wtDgbkZtZFmr1yLJz0jij
Dlz5+8KeqQChC08UiFWy2sJ2oTo9PBLSYiXfT/B3ZposIu+9XlNUx+w03+7KzGU/5ltpw6+GnXIj
d9ewL9bf9im9Bs0P01Yuzdr8cGOOoqB7zd4ud06QDLw/vD8BQQvSr8yjDjYrqk5GqiTuxFN47EJv
n3EU++kl3VHyPl2USrGUW1PxH9LfzHH9kdwwRrE92TfzI2rcPdzRw57i05c/tpB9YiKSHTfyZBMV
qrrHfh9WOm7HBUU1JUBGshAsN1b62gjjdXDDvXF9OiF6cu9JfT9f4GEVxFP2FICHoGtvR1+/Ly9w
oP8TXKhk4FtVkdwnIL/2lxECB5iUejtJdXYLOZOjQNTpNe9FnTUKrt1z7sFT3EOuO3KPuanLk3Im
psUd2UJ6Mj7iOc3yFdbzUCBHbSnPhztiYEf5rO4iugY7NRQ9wq+RdeH8OkNuS90G2C8zNe/fIRni
cCjyEpfs8NF1J78mWta4UnH6sSyIrIfIxzAfzJEwlCndvQo6AaGJSkGlIdH+vlQDZ0Pg9WOhqTgh
F1i9ZEx776uSpG46nbV3j8yGAJsb7dsQdr+J3pmMU+C5/dd3JkLewEXX1CQmanN7CO/xIP3YmiD9
zb9RQtHSqqmiRoetSCD95pYXD/VVl5j+FWW8id2S67CL+wCQj5sJO+eKSxKTIs6dQKc7RZVUyxDL
iEo8jSJtRTjCh4gM1YdK2E9jf2eRnoPOQgwEi0GtKZ9j+6x/DbqwGivJHt3KoOrI9AldnDBWi6tl
BUY+IGvfMto2VRDxfjcihsRUyk0uyUOKpLIuX4fiaoUBhbEtwbKzTLUmGslaHPiBfLm4k6Ff68vd
bzJMF77pdYfJ9wa9TppeepVMRb3S940CbtaCDDnD/l4O5WlwurjRXlVNUsb+/4s1BEftEE72an3h
WZ7yVWzeO1Ts7W6g8iv2yzZzBShP/IdWnerWeqZ/NeGL+hJZKntrTTsCXeKdpvOIBHOQEIDfp9LQ
zRSRHpSkWBu2ulpTFNZlOtzruU0fRideavgkE3wUdVFFFAFdYP7HUdAKGMsgGUoBFWob5yfQsHEo
YME+wKV41W8VYn59DxhG+a/j5rBk9lhtgKkDNiZibypSxs0gGjCFYuQmg+1Mnlp3dwn3py7uNhEA
akGeSAQnzsl5IOa3NVwf5CNjr1jEZ7pvteG+iAZNRad4uPkqls8i++CMEwWioH0ULqXXhY6xbo1j
gdZMPgRnVNnbSVBWlUmis5RzDAVY9qslxhIwiqBZ6JW65XIZvt+WhDJ8qcRUcAMUMvzhmav7ACGg
+2UMZAp/r26mPnA4KmOo3yIXb+wWQBaGN6zPo103mCtHXtZKSjcivU11mZPKgFgZGfTKlexKMqBb
Yu+Y8/ocQIi5xRASkMlt+RrXaLi2a8OUwy7cMPao/sJyrI2MIaKOa/ns2H+3nM5vfekXBs8H6fPA
YeaRDiZfpfHDbuelmb2zQadzBjvcseE8bmRMjW19R9ClJY6ZKceZwvgXtvSNzR/zObD2Mk/EAlLT
F/sfSk3q51PnuaDtMMaslibuAcAOdM2VgTvYIHaa9iAjUufxZl2teC7T72rmBw8EK84DqNKa9oZH
+RYssgExmNT+bycF2mw730ItUMSUPiy9xTFcgLGJA5D10jDnFLYwmU/ZeMJ2x1V8fQD5oK2G31oy
V6ebGRaXrq9t3v1BWuKCYohGckhuHlaGJTdz1YDLyTahsEsfGnfP/+zXKKg/FSHqNmK6VlFCwEWg
fdo2YRDj8bY6ZYPrbDmedMfhbaWyLrH6Wv/SN7eWXvuUAMGXEZEWcZiRz28eBAr3J6sW2Gx2tpBg
gYIZI5AwHC3Rrf1hIzBNQLYF2WDKwYZAf5CCyZdFS/HW86M0RiG8VSHINX7fZHfp8dBcgjgkd+KB
PaSZ5IWQhS6+JPD/CTQR3nrxTHG4BrJ78FbLFqCY+KeJkZxOCm6tdIoG9ABx8svkATs/R3nmkdW3
WoqEJ/l2MAO27rCwk5hHV8OFpmd2WlSUHq2lhRpGlHMX6DU+HgfXD6EmrHxqr11odV82tszour+P
1ebFriNV9x2jK2M5FRkVw+mXnxZiz/sbqNhbEOOUxKjCTZKA/L7m+CMqeayCXHx5GuPVc1svDviW
ItEnz/EXU7NK8glV1V6qcketcaGPCfii6Iwc2nDnwqGTMI8nL+ATCqA/2ajwRgwAjKUIuxF6C91q
FV5WrwezeOEF2bfBDqVFOBQBGeTHEu2/8gVKcQE4Kp2YIV3A/GxySC9bqvE1VtwLDERM4nhcnLdm
Nk/zDvFQCl3R40FdigeACr5c44GW1VdiffyrVSLcty40JJ6rkEq9MsnruCEqzDKYAacQ5GtPqznP
vL9qOtXvPc/cDyaWHOa/SC2r883Rmildx9iwL68R5qjye1Kh07FW8IoViHc4zBcAiBoyXiNsrv7c
+7nCmErOhB++lm2qhPx/SjeU2qXyMabUGCPCITtw/FlHQnO6i1isfcHJtjskpxe+3aAR2U1XSxTu
YKrhgdiwYhe7hyYo9Hqys8nS1MfjavtcjM2Z1NIARx5hsYLIjbyD8VM4q8qeFAZUUNRR+22bXy+2
d4XtJSrkWYtdj8DvP8XnfMfqhcj/ifW7qKQANXrVhanMkTW9VSm+U4XzifGIIKqXGgPsNACsIGLX
43P/bwKbtZNW2vHgI2wh87rtIsafSYe1MWOhpZOM/FD2YXa5Hf80DYAD6f7A1GS1+YmsAgXRoD1o
AR8yZVO84uGfu8v+Zo/ys4hKCxjIWJwP566dEJxY8yZE0DcUep7ye4hh4cRi/v4Xhhlr0yhYaXk+
C+427nPmuDClG/Od72zbwJ3wBMBYpyped1eCh4AgXCag01D2YukK2lsYoRGz6ipPgX5lQd5xO2Oc
v14uFGOLkAZWnTD7ElMrnHs0SD1wi5RaC5QiiJ7/3L2bj9v/alkH0/yf/q4+h2iTUlod5lyCu5uv
AEKalW9JLD0ZcgNihTdB0AmNncZOAcn8gA7gFT7gAPU/v5KUtm9psBPn1J5MAMip5mdy40KvyosY
kcoNjXw52urCBY7cv1+weJ3rxPILOjyJnIq4xhpzVkCjyJCb2DXsj+92TCnjAm7WdMk9rjRu1arr
zuSWfH2kahAZZd2OZaTtTB11mfD2ZUFrfptukkwmrCwtJMsJDSxLZFgYGyYamzRZloIrLa8Adoy5
f7kiRpefWHXlnGlyr2W4c+J44JPZDh+VAkViQ36axwuueuWcWmtaaSYjVxWJF+/yunAsxyZOsu9B
FiMTibo5QiFZ7r/wFN88G4FDA/bqm2tbak4u3L8FYGe2t0qRrJUa9alv1FL8PO32HaL2JwRqkAmV
cF4MOOKrxeCEpv6obLt3PFHAYE9oTwiGrDGL/sB206C1dTCzofbntNNhAOY+MocwqWbRxGhyrj94
Kpbyama+y/OMhOGB5hC7fcK5Hrte1UYNYdv+da6grqqzt6tSLbaR72xdI7zLbXq+Ekqt2xK4mi/z
hc88oh9huJEJemrRf7vMq7waQKHRBotbDKfbpE/uwSpy8N+qNrM7FepboxapiO5QeayX+5yKND1b
6m0ZqfoEJ3vXwSNDOabJPq8my3tmeqm9dWhbpSGzeVrUfaLDoRa3gSclhg2Hxg8mZvBdVhgQ7Ic1
ObNQOgNju2PXPvuvRo1uNl7ys/i04PLOvsveq3W+t8VP9fbRuGitRjig/YG7VabUbcOcStELt3MP
BZJ9tP/EOmHOgRDb3u4oIU9aj7wVSQOpa81+3M4y9XudYCDcGxz6kuM58YTFaAigszNRk/5VvA7L
a70dUfAq927xBWeenItoOLo31n3tLJRJ31wPQCRVdI1MEfay7eBxuh8zfHHRoIDDOfmIZ3yTU2Zm
g9+pGmQUEKAIV9b6Fi5SIOLLrCu6VAfkuMVCra9ROAphKfBjab+ElZtl/X3jRz0KyuOBWR/mZEx1
wMrXyXNdGsESGSlto0ZyhzeWP/n9h3f9WkKl6a48y9QLcwBsG3GieGAxN6Wea6vAUqd/Vlyi+W14
raGNLYjHhpQuxc681emHT7WLGRFzZ2RHKtCfENRe4Jm70uYVCoQZL5PcKicE12TT+tgfRpuJ6E9K
mrG+nrhVh3f/48P9ZsSNg2A0mqzZTzPLONN2tLi/T0521Hmlu1S1Vevrr91GErRYiHOa+2T/yyi2
aUq8woixerkkPqcqwrftHBgQjKy3NqYnrFyY+3t4DlPh2yCC5fRYjpugf6um89PWX2cnau856I0I
mJ+JZilMdKdZso1oXvHlLVdhEXkFf8s+HEly9zYwtpepHX1m8FFTBejxVdvdwI6C/Jdn1Hqp43gU
9TIP7bhR//TdJr2MaXp5XVZ3O5R7qmUKDdh+KMKIhHlslfP9JDmgAhypV21a1hgkKvU6BHjpqluP
4K8D4Z+o+0ED0meY3pxul1M2dDxPlFimKaCAG5/qSdLq43zQLYuyrU67KI0TGWQh3tiE6xSc7mVY
2ZoFm/eHZJzQ1psVPD3honszrFnYwlppiDcKJjvtdN5XJh8V9slIb7dOuO894k7GiMcD++DeeWhV
fztUYYSxDHHhPhjtr5FG6cUq6hr5iHj/NyvcN7+Ut8ZdwyVeErbfuAgYyh7MLBo57mDwXK/JrXCz
P8ckFdT9NS5LSDE7ycvFFtW7+LhiGnSEtLadQ7Sn2h0DzKQqXAq/2BTbZoiHqVdVhWMmV+Ykd3FN
CkCbF4MnTnIoU56lIbwNkpnLSGT1b95gwULAwppx/S8OPOLFkold/cE36PnTaNutTqppXIiZOvfh
6xDkugcT6RiAiBzk0Ph80qFSvnC3v1YtSNFU3eghp8k1EHjKXAUgH5lcO3YGu1CNhZI+9B5QG4wx
86zRk8VsymdXZtdDF3HV4Ybcq0RcAm5CCW2AMdVh7CdveT57q0pfv+XlZVj16XwzuptA2ObCESpp
4dl7Xz+mU6ohQhpZ7fGc6Y6vD3/rVEN8HtOw2+sWPjpxAFrd3OK8Ef4I87tdhcBwM2D5NEyDCiow
OMuWbIlU2CNg0O1DAY+mZPl8IJFHegN7bDDmzwjj9ey2f7ETCowkFRtsCCVnmkhlFsYaP4xxCVlI
p72WT+AtStCHnDiKvKkPzOWQBYgSuIAix2D5HoPcyQkbqjDU1+r6YDhpCJk6dCES9Mcew0yfhOS6
nVZC4+zr41x5kTcdyw81KPZr9pXkpWfxuuDV0TD9ayohgiBkz29HE/Gr1iku7mUIiSY+UsVASmgW
TSPOJwzc7YoWBmr9zOacHOhxOT1wptGuslF7pmlM+DlNj1lhwQ4lUTywyCrhT5FBf4ezOfNzjxkH
jrwh2fMCqMHWuQxgbIwHWMlWr7tgIQgKof44bjB81N0w5bIvDfYY7E70RjruxAOdKXvYrjtamkj3
m+HXMkbjamgOBF/c54kiFfJMGC75FUqn2fjmEbUObSG1IwpP0hb2LABejb4/XXtUCegfzCZEohtP
/ZrQdXDKfg6gzZFSVW/zOkZSs6MPltyOwMBIMFmBwxPSqoEZatVBmbpIaBHgw04iF7atu0F1fpEv
hMjejwQSQCUx3IPDj1z2U8GjGRrlbyDpKZlajOg3SWmH3Ota+cPmlRPvy7CkZ0htDPYiKMoBOv7q
loQ+xQ9/1WHI0poWD0HJvEHHkSkFY0Z+FbRcxcUqrvMs1uYONwJr46JC0kBZiLrOUiipzokHuBF2
f/RTurbyGzWlvUoQTbjB1jmCpK+Jg0Kc3Pjlvuu2u1FGke3P3xFmgReqn4TKbioBvDoC7J7YnTab
UM/wPSeF90KOzrsXCtAWbAU+AmZhlNrOGgYYIlc5g1ALd3ggRSJdLpSJ7tD8HHOkxcsjZetuuL9p
INNcwtzbfmbogkL3v9yYv0ZGMCimArMMU1f4Xy2A3Rs7t8lCwEEAJojFaSG7d0qWGMmX5R8ARP2+
Lz0Z4tY0WY+UuOC65NwFU1kmeJAiFLAZHjkcBlzFaWi5Yl22WExhV8t+rVOpN/aXJwkXFY8kZ9lU
Owy1pCOe/xz14cwuXHGyq27Js1M3tvuUYtBzwkqH6Atf7ARfIkMzzVFiKFk+2NDl7OXxLhNPIJGd
dySxgwy/dga+vANwbUmylvU5lxpFaa/c2TMEp2DzRd1KOovORwtjYOHB7M/r3hsFr21RDDOruKn/
8bjf6rwM5AWxjAhnF9MB+e1FDhVw2ic/bH4MOHm95/6bUMshFLBhUZDd8suV6NOXxqimFwIYuTzI
AlfmU8rC8whRUPg7v+9UOwIYSEnlzRNx227Cxm2ZDNbLC+21lndThAC0n/3quakBNpwgE4yrDqef
E39ynAQgnSyvZ8rTyGSFMc1bqzTf4rGncnMNnQdYsMCppUBLsfQqQG1yIRR8U5olTIZwnw9Fe6CN
KG7VR+CKUKlY+dEbY3w4CC0Qx9J9K/T2RjynZXmlnJRKQj2sHNKUBntfmJRNfKT3xvHHHuxrOss/
7ZSmMhDHVjz6xSjLOzlGWpRFA6lyFxvXBp0xLM/nZ+w61vMYpkqFePWq0dix/GJ05RKFsYRIkPeH
6K+LQZuoO9xx/pRWt0445zg5J+1tP+5yH20FIBd4uVJH8eanpe14s/sVbNq/4ODEo83wgyzq9tK+
VuKcHZHVm8Ks9vAz4pqTl69+USPj3VLEZ76JsAiO9AOUm5lM4KOT1O34Vr2mDKn8lZ20GDgIpaBm
8i1uq/qBLoq2oKP9FVLA/c5NwxJo0iBWbQrspwKO4Au4G+V/skLSXv7srLU1jiyKrgo9j2ttzM97
glWNdT10To7tHXT9uAlFRic5EtyiRwiAnxtQNArS9nk4zUfLzaCfIPIHi7LJF0h1SOlj1SRTxBmw
q7/fDVLZ80fKSlGwUBiV4CDSEGICwudHcwN3DRZhKywyYUOqJOkvsvUMjnv4lKIir/OMJYdZn2UB
CbVmDwpqY8gp2jLni1JqeqDEMzu4Ns//F4Hc0HEMBSJyamzww0k6K3z1SkM4ytDBqTHC76Pm3CPc
uQ5MsztDWfptikGk5RYFrUvhhwSKZeMIWmvt/SGH+4TrFSpx1PM3RVZ1/DDEBgxKaQ0UoIwSH5W/
bt/VWD7xgYPAJ76KDQTFc2TOGqb42cKOZDjtb7I0qXXOpPVweadMlt3hYKBVgayDW/H6dzNNmbbN
i6HYJ7UK3X1LSugcWjfDj0PINvIZVuw6/DyPDOsjNeay/59eo8zb4BTlVHFFJVQ1ACeIyX11Kajp
WfLCHkyYgSUx4OEkmL4cEW5jAnSye+FP/w7m5t+ym+8U/mXv5ErQR3w8JVgX7NbTEmB4J79VNbZt
WX4wY6P48WkzVB1GC7aoVkfhhaz3M6VkXgQV9MNJvRA6sPwqyw6T73gdJlAmd3yCTYedKkVZDuNn
+fRTYp+eZqfS1qugcRuPu8aTeQpHxhuOWf4GuhCbl03/y4+IPoxMOEvVKcz4ZZj/nVEaboXTDM93
VGc61wU2YCR6M6OYQe/na+rtZeMU7ZMw1mdx8mRtIJhTz3PYNUIufSi/EZax4/LxNepjj6mmHVzd
w4zBjMV2opHpeUz5LjRJ9tH++JcfyNda9kYsL/sGUKzVWLfbMciUcqPwrTmc7PWGVc4KKhf0YIdz
s4A/VNyZw6gVIlfgT9fz3Ap9oZ2u5GFCjB5VA8leDaMwjMhA+It/VmrRhhv6tOp7V7OMeAm3lIMw
S83W4DwExkP13oJyIUakuyOt8bt1JDnmP3XTexnDR2IBnZF9qDuTa2ikd0avDDvPvu8Q/pjx3OjL
fe91LKab+uzMqaLPhBrz9f/35aA7oN++3NtU2eAPN3RGZfOQaLGwxvIUomBjsynXFd2MK3DfTuga
XbvWBn93wMTAkI7yZkMTdsJjT3raLrGHcJ3G8jYhygM3iu56XSZiF5LuEvjiJv5CrjhSQ8FT2DsU
Wmp9QaezYzLefA7t+uQNfITpS50ub1nzc4JQ62NytRrET80QIx/KxMx7uU93VyeIPlHe6FDsfIMq
nuLwCPY6FUUdCnWcaM43u+wE+kNBdb+jiyVKBti1RrAAOP/Hw62JpTWe+A2v0oM3qZWfN2lSNkXm
fVys6F1BT6pwZTYan8ugEiOEf1eBXqGhYsI9II8NPJpkEFRQe79jqpOhsX13uF22tybdOuJfl6ql
m9sYqkmX1Br/PXVS1Q9Q16PIiU+KnUXLkObxeC+WmY6d52ZRaX3JsIUoVvSEzbxGu4zslgQ7I2db
bhCt8UT6y8szogNKBHhItJymrzD5OsWXhJSR4nga5Kb0GVZmwyYFlqjUfcm353J6caxpDtgxQpBq
PzEwkkE3Gw2LXpsLO0qGokRBmgiPeGfz11PG0GRn30N+Gu65dbUCpqQdvqQs9vL3KUIANwzBH4T6
SMn5l+KBHpOwASRWm3eauM1airRWK2wU/89aKetAgbPKUBU2J221TdxFdcViTgb98oP8xz50/zbX
2go+dLUtODxxei3uFbplPwIWfXasw2ktqm1YSWbkGUmYbL62L1nMxwVraRP+hsFG6n1KrseYyfxa
u9q704xLG0O28Jhrt//OnbDTRyr9MH4TePxTOfm3hBZrgC2NLgpXG0gSoLHQlkAFXIlm0FOlQGKX
jbISB+Dqfx4CXRq1YRPx1cd0BTnf6ktvIhWhT/w7xxC7hxRJY/bws2BK9eIEEuOsXLLwdYaQ3M6P
Z1kmL1V5lMmRqPjYRQo5lm/qSAKJ4hKTj5hjyY8sNGHeFC9zLal+ET9mFF2CkzWmQtOSGDxkd2AC
DO+paYwqDw634Ey5vQkEdvygCPVmmmpU2Jfhu8Z53Ewu8oNN0uIL2j23z81H+gYnGSnXWVfr27Z7
nz3cPIYMN/FYLkT7OqOBB3DsNL7yw8SgDNJjzI86eGRBK+DEMBtEe9pnkXdHkXw4HMG05yFUmBey
HoNDDJMXyLO7msCi0zjZpfeccvkPs5Rly+fX46xRCyPdPoRINPAjBe4XQLHUIjIiILxz8s4AMe1u
hx7IYp5ED+g/Q8Pkg98qK7g02WOzjFO1mIVhRnx0tTps8iiaLJhGi9+uCOt5A7vtCFH2vwvD3Ad/
LaBTlELyg1314LjoDZSStAaMpkMOoPEUFCS3EU0npO8hblpSSWCpgagJsgpGYXHL3pekQYBgByR+
eSzASuctcZ/oa1G7cBOnyXj/FZ2BUIttW5UteR3AgrddIKS0AX3WgTSrXg5LINYw6HMI8jOqbq0h
warqlkOLbQSAk82ZyJZqChCn2duOSZmBf1XdTfLGUDIMV6chm5Lil00CbnJ1XWaW3pgiP636TWiM
m9nHI8bCub2ZuinAIaZY2CBXqDRdH+V8CTBN2yTF1QCCZpDDW3w/n+16LtTZNDnd//t0pR3gk2Qr
/AujD7YvNL6s/oJuI88NRv7AC9vH+e4aeKgsivxZXC591nQCpyXcnKWcFgL3wmwS9xE7+qtYF1Bd
CMk+xgr+ykHemrJP0iGmnMff49fOLAVjQrU5P6Rv/Gq/S4WihxkUiQrt7Aa9DFIubVirISQotQaL
oPkfIrXdJrFyZFmee0Z69Zq9+ggwBBs3q7XbU7HuYiS19OLn2jYS177SiBbOnclkYrFxBMzykYdj
iu2L4U2GpHOrtJXE6OFLpcVzfgAyJogDyX8U4w8Li1rL/xBXvP9g2EdaPbeEk5Y8cdDKwacLQ58v
fwNTExvBRNst8uZiyKotpdtxQSzlPytpX+W5KPtr30r9HOrNbCNQtIl1Vgg2iYesahEZ6CXUAtDb
cTOquR65KJs4tSbM52ScSIyF+GGmronsGn4gbKJvl2w6lQ/H2qlFwQxK3jG8m8Pwep2pdQTImO5v
H92rW8f+iATHw841pB1LuVSFSBhvgUqn37I2GXdeJZS/ceWqc+6LnZYgpEUhUzJEXnAyeWQVJa13
gtv2dPVV9aLJqhFDvVfPWl52ePcrQqFO+eD4z5ma5bxns2uYnsyK97K7O/uqZ0+KsUrsFTccLTjN
jEMs5iQpqb1ZHd/m2d4AB03ItoHuz88U6p2geoOELKMyDhZPKnzXmpizF7bzyvs5SbvWQRWr6zG1
zpjJ5G6nff/iduvvVxz/pITmfy82xDKwr+2TL20r4UsNkZ8Sjfn5TkedXUSiBsnxo4mskGo4T2el
OqfBIE28WXaxx3Xpe7F99jcZ11fNPcnNCg6s7lmQS373nmJFHXfOsASIqnrcI0YuV6k+uoSrI0e+
N+oy2YbhszP/s1NUEgCZ+dVBtvtNyaHke6a3b+7T3TB3bgDQ/jbtS1WyZKYKOMi2MJ/QpQlF9DvC
RzJZnKHdIdUWlkB73beO/Q4A0YZiTxNRNaIR10dSUe3HelzaWFe8w4zwowRlIEN42K+ZNCXnVUOb
UCoXN2fN+HBNt4gIi42pPGBhCvP8J3qFPsAGtS/8pVRxVYrr9WbwySyvjKZOiR06R1/tTRjDRz6F
crVoWVCKJUFPJyl4mGW8liUusUoCdIo4qBgkWRjyO9SLhHxZfvijXEt1iIldqD3zOFZkOWvezocV
9m00jZ4DZ+B3kgAssoSkXjPcZBHxbXsOTI29/VhDKSmXjglxtMDYMx760WP+wmf+1Ul32IhnCcoW
NFCfS+vF5LP0GQ9ATXOiM0Ki/NBIrhZ5rj+oaSaTAW8wYX0TJvbrllkT2O1+2ZIy2k5WbPPn4gdQ
xestfAmogKv+1RZDdXIyioCxFFaSIxOyoGLiSdopo5ADL0mYTQVe7nZS9ISHT4wn8o1WLCr85DLL
TER4R//OgkYLoTakU3+MShykC49mvOyXYpMqqskTmKNZfNBAzTcpIFhVL3cZDkbIoXhdqzTs/83I
H5Q7qoRNihhoY69KAaFqozO7AfYsT+ZnQUkP1DOo/CzHbk76/wF9gdHtyZl1dfp0p34gULmSlht9
LFCY5xTmEyE778mr6EhEhgal0EovO3XqNDyv6UYufzt1lunpHlnkSCyhu+37BUV3CS7Wz6CmBKt4
SRtC4M9vZUqyBUwE2PSxICEQzsRKP+NF13zn89Wel8Bf+9mEtPSNQuM98Hd+hUNPOLPhkl1iVYMq
G7+XioxG4pgS9EHhBku37zeijSmYWNR8zMcsNGGBY9iE+cux3xfk3HYDhhzoMhzRl66JaIAQ4wQ5
ohVZMZSQu5Kqc8T1SwLF0arTDPWHu45Kg7jTPJH31jxbVtk7N3p6WkOrXf94R4l7q8ZKn7B5/5Ch
ESggB4Twp4kGR6Hc6A0hY5v4D2pHc/pv7O1AHUpsxwRIhY/kZ83iaXLrIhDSe/Zphh9G4440Z2bE
z+u1bKpUSfLF1teoe46jFEd9KVs23SUuCHrKXOqamXMMTGv1wJqNn76BxGv6RKTBD2DxwoIXRtwT
Ly4p5XFyTz4vtM9+zdL0IdWd0I6PT7X20P36Hi7UUyUNAEmKIm7ECzVxvI9TWUmJaO5BTOYOU2EI
bpb6A4d/ND4QbmDwvZ33tn8SHRoD6ygKksuwxMP/MOUiEPWLneEBWhw9JchTC7Ss0Ctiq/XBc56Y
33ehHpiv2T+oH9x1HOxEFa5VzH4enTcn4v6U7zKxR/QIxlvtgJhxPq6ucUGvfnnct9r3+X5qCqEA
CrFOEzHMOy1MtSldgQlx1bTKFhkPub/igzAG2dM34nkWM/k6O+wa3LhRxmKF1tvFCKcqFg9KuNmk
Cih9pV1Dn9yrdd55G2ND3YTRT0H8+faA3K+79dpFrgEQVseTyJ/rcf7P7g5kQFIhOSFC2V8/nPJB
Tiz/LbiZSuD8DDtfPDm3WBMtf1EdLxsB2HTPGmCwBz7E42N1e9CG66gsOgP8ZedRPEjTxva/6lPG
gQg5XAebUtz10HmwUO5/t55H+nB2mrXS/WlyqhJ1pjSSpGCjsQ6BhuDS7Mh2KhPIR47b4XiQDCOB
sQVwSFZwaSmoVXcUZJn0g1jQgCvIAPUL06le/YfYbB+729y2COjwSASgRw2wiFwaL4DhoXLEfmJ2
aenUjRkh9RRA6z6arFSUVkvggEQfx7BEde3wfk6Boij8UmhwybRo0EmhW3lZYu/w4RaiVHDoPdm7
1z8hqFiKf6dpR2wCwSM8UdrLT/HJ2Ah6CgSqtXacbCGeoud3qPca0HzlbKWJqKCqPm/W6ZhjNl4r
sR8/ogFHNMfR/hniEy+9O6FsWGoeR+mMPxpYVHHewztlWfi7IG6wlS79lVuebUrwoLMtM2uiiz7P
ehxfVxk0TM/3jWmgNpKCmCp6atpL0cQR7bLsJhaIcOeSBSvHYQ8idKAnRwUjvk2KssObBcY3yL7B
cPDkQFgck1WGCdHeXTRNlv5GK7txL4CZcppZWfvk5mZKyr20mKTGhJZ4ZCbKdBwTATwyb3axF+td
iSuMGrK4kzXJlJtIRbDOAu35a7CY+E/EplgEHc6jWaDqFrxAricYg8vzD40+scvWcd7QSKN7Mt4J
L21JWPnu2GqV+MDsyndxLRyC/wypB4LrOgln1Q1ch0ps4KT1tJtY1lhiFTuL0KyMUlCTzax/AqWW
Mgv4niRqSJpFrVPtwZoHjjEeZATS3UARid3D5ywpl4gAyCxewIGODKvpbmM5twYiD3OQQvlXmhFQ
U+cKzSxzU5CxLSpM/oAlDFEE0N2rp14Lc+w4AM1wVYAzzFKbdaDABNEcfNP6Obd9buH63D6baW22
XYHAsVIxpp9LNOi2dZQ8bX1ZnU9HNyplz7/P4amMYWDNEppY93tkVEqppfjbQ4E2SDd64CKg1BRK
yrZOvdKAqYoVbK2cvnXBC1I0n/og9Qsf4eWwL7XNA9WQDG0pcs2OZubxKZFaJbFUxbQ11ORfwA/Z
j0pvSIP9FW/hYwjIPQTamPHfjYFjYoRCxk63NiHUghMhGw9X/j8BeileuW78l/uBhnYBFNvIvJvf
r14ZsGq2k9aOPAxYISIJp8aMz1CU+wmmE8Xg6OhkNGOrGPXVeOuPy085pUaxBSQSyKbXYlzB7eHW
GKOy2Q+/+cEXZuEU3QN2DXHTHp2Se5gDrwfoO50VFhmBq3RqAwPSEYBtPzJdgkOdLINUf5hGBzJK
4wXVF4t2T+117ifh+uL76pzbTWXPMjJmFMspxwdKaHfLK9YWIcbY/kNQtsHU6YX9HKBvkxJW4PJm
wLP4M6dLSMZQDzbt3i4eJpDPNaOA1FGeYIkV0Z+CEDyPgKTH9I285aULPY9hmAQOYmwzRFQp4TOB
EWIVjta/2XCxuUjdVSRtMdBlTLHVM+yePLgaWqyhTVqx/+VKu0K4kAOSC0TYVOPB9wHwbC77FksJ
5+zvqQcHOXIS1b9QrmFgcfess8ug5RLbCwS0lVmlMJ/vP0J5/2qRLPxijb7v0ernliaFKJ2YOdes
D6P5q7EzoIkIx9YRI6ZvXQxB7fpIslmCBZsqljzsGX97IugVJLd4gzCG4YM2iCx9e4s19eE4oTFa
1pusO8lYUQu/OKYhGEiizPeF17sfDR3jztB7Joi5sfzekjCE4X0nF/0YgEQ6jOr0cFnXIY17or4+
3q1VjZpBrUBEFNom6W2thc1/At6ZJRajBnOY/cQFlQvgFPkxl1UsCv8RgO70JaI056aagWWn6ePw
0+3/2RaEo1JlG7jzG0aXbH+gL7yK+V7F9ZA7isvphI3JhDjKdN9NFNJ4EzWDa0vHfHlXLsGbCGrG
QN6ficMQR+kJMibktna8W+rAZNzrcFOktKs30FzNbzAqahpdmJOOG5YHKM90EgG0HZ2RyWWZ9XHK
Lxe5uj1/ptKwjN7o/JngpnppUpB/xeAmsqMx+AjnhPPdcumv8+XSQ3/7V7ttUot3YMp/X1VrNXjJ
KUYoRDqms8on6+8e3NUETFemqj66/Anedfv+3DJcky0yTn1ewifyF8gsoo4WZIC8kXheMHwoxdKd
ZrpBvtBn9VCxHSgXAy/bs0TTKmk/QPqosA/yHHTL2rSJlnxA5W671FGug3LWaqLEJij66YDv2M73
9YNcJWX33rLwAqAe+B1asKUij9AVzl8XMwTpYQfwhgUAe2oKrNAYE/FhAyfbSo5qVOK8pvtrupIk
infnzc1VGDVNMvM0MYYtNnuluDNLSbib/Tjf6qfZdhGUag8ySU6+jkZY4yINBrfLqZXoV/WK1zxf
gBAfW37hO3RAYzxlyGBScU/LtOWmJiSFTo1Dfhaff5/KGR4oOv37FpQ9AXnU5IyN6jLIdbWIWvR+
YyWAXsItFZwQ0ivyW2eD489HyjJkvvDCSX4lQOWJKaTaE7C15iY6LLvPkY5mrs6d87KdefzxK0j0
2fpPmFM1l8K/ZilLAMs9Her/IMV+mjyZmLsMoD8aHkbgiuif9fGnkej80aWv8tuI1RGxG6F+4eS9
2+xuFxxnhLZOA1BYinB1irp4LZoRxY1jG0RSsFB3TPJN7sr3Ang/QKI9OYxLQ/eXQZr0SnNahuvd
niA0viTep0RCz50J/uj8tE0PtqpxEM1egPLeqTZNcH6xWhYj3btn4SKmY5mGIiJyikxuEZJzDCrG
bGthZT7TShcVNnxTKqNKJHv6n2764Jl3zR3WK2CUELrxhZNv2cs18YYOZyNoXi1Stv2ZstCOCSQU
ugTxjwFl9ykyJjsgHIrw/SFFwq/0pQdvvpeZKq6qu4x2KVc6QJZEFRgchzTd+WRMPQutArDpLegy
CdvpdictenuLOgra9JR3oWma30SvoiCrcSjP+eEMW/YMg/pL9mHViXTPN3MyQGQiDMembGm2n0aO
rurcJDAUv5puCV2/+kDMSCACgm1TBcSYl3eInsULi0CjbKrBbg7CTT9g3oE3TluxTbr/Eqv5wAnM
KXgzmNctDz/V3l+GXNNFUIIe7WlgNT/ZsvSOO4Xm+rbnMTXLJhZHwSEqmxx5vWZVXwx/S7XSGGEQ
IKkSMsnsH8MBPXbq5d4CGE4IPbPDwvWZyzvUFELF87aRuKWysaDz9r2Dez530mhTdZkVyRj6Cnnh
r3c2Z1y4g1zyC3a89inlJw8L32QBqn96VtMvcdTTC7PRAURFRtb+tsnc+j2qX43lDF5kAUqkDSsU
Q22Eh4OGDGKxIYa6nMU99D9btqWJWYgV3OL8s2G/O0i0l5ca14kIb0L1ztttjFbA66/gAA8J/TbQ
4dppofVy/nYrZi6seMjLT/KEFJ400D1yfqOtm0wCeTAIa+NuhoJEVfpNQ+qEqjapYKcuo+EgrUmh
cUr/e5AQrXjwkSqWz8eaZFTmlXwBfZB+z7o8Rb9SudidEMEA9R9W+6Vfe8KbA8oXo7WKdZv9wklc
3beExVcSmkGYLJsjuq+I7w+Is3jdTyDouIlE7mecHha2wlJJrvbnmNxclhHtGVxkDJuTwqXvIDPP
2AenjG6RsFg5108/mH5mJUZJ56wQx1mlwiRBXY3ADLo98+cQjzyLuOw/yyDthNmtCtPI1qiJtW4f
w5VtuRXkEHw9OcZjQJfHSPlWJY8PA4z1E5BtpkYsm8InHyQupteJyGVbzuGMlXdcKkoJE0HSqTnq
pnkti8snWIFhdNKx9O1RU4Es3MyvhQbK5Vvli6wl4k5sldbuVWCa/en585giu93oUf/D5k47GyON
ZJ6jAB4WVEI78taW3bG1qSHYCn6KPMsF1lqsJylDXzN2jozWbSla1nD1I4dt0jTj5XZSqtVkCPSB
ldk81oTVHHv45meQg57C24O93dSj+b+7QIxQwdKSOMpAR9CRtLpUfWug7FUihxfxULvyzI4Yhnxj
SgTbcsXdyrmGSJNAbsTrzlJxxT7KW/4Stslvi694V4sDbJ05NwEH8WZKL3NCOA+cxdLuKTR8oUig
8rm9y1CN7jAXaV/RUJvlHSgY0ljXZDshlzp9M07w2WDCtlMJhuUJ2lwd5nFH/2aCQAZZ0nX+16SS
+/bYJu/TqHxJDzc0RFV2418fhuMAZzO5U2DYhKdR5tXdomcAAAVrhSOV+I/uQMfCV9nWmL+Oq2aZ
Cywkvi07yS+kORNydJYANP62f2/D+aRS2p94KTdOEzW83/DXDZ3feSJGtXYf8R4gUjun36QEZFSZ
fEwiEF0jd1qH3Qsrl5uvTjU71bJt7bZamidbWDczoVz53Xp2T5QqGJHPHwwFymsHzkiVDSTyC5Cm
lQdikLJMXD7cA5U3YSOsA8HtQcN2PfZ9h617eaZNZN76DVNeDBs+9P5p27cwZDg+8dvyz1jRiwZE
zKLysLLd2cQpm2g1XUBRXgakSboVIVO2v5ea2bUFU3khioM5aabjmU6Y48o+d4aXDxgDf7qJfprH
fkuxqlDLYUCqnYGfiKFfEhjn4V46IzqqR94lybcrz/jc9XImUvPanDWWIRpuJiJehJLlD2cxbfqJ
9cIXD9qbcO5pGvQxyv8dOQYhmXRM3O4tbzhI939cG077bCpRs+vOM0eXkP/yyX/PJwpCyqVH0fBQ
ZxAtfML4fidMiMrpsyQ3mlJau4Qmc6eMLJF0qDBOZGIZRQ+qQE8DqR118fZkO1FH8MmvuhQy9M0F
iCtqi6SR7Wuek7ttV25sfGukJ62o44Scw845aryrbBqVhkBGVyDcL35Ak5Y6KlU8f1B/ionkwWWy
aMOLvt2hbD9nhmGhVoXtIeZKI9fcxVi1VDdtnmDuN91nXoN4ZItxhvVIcZL7pkD5wMr1vsBclz0B
90jUmzZAFf2Jp0FJzmmvVw3YkiNUwZjS7r6iz7C28q+2+eyH7vHqlg7JFirg+z9itSqfSzO8fED4
1nzyBTtZq8LTdF9qfXQ8gioaJZMWjovVgNa2XKNHHsAe0S2Ga4LAlYQz2fK6mLO9Ctckq4JulD0+
HHmviZ8Ee8brEti3CTXTRQod6oCO12dd+EjfcgkXoWUhyOrO2dvUnZO4DSGtgJGsrM1XAGfyfnoc
qTVQgBX1aODinF+Z4/kCWeaUPe9bpfwxsnrCfB1nNXcTCps1FYl6k6IouxDYZef+JBis1/uLQAJ9
lSROQExG3OkSLHKvpk/oeCKzgwyDjiRpyyQWibnXKXLqs7bMaPv+uQnJndsQ9NVNuac8il+2WNpw
I8CiyGrskDKalRQ+pdprRTzwX1UmKY5fjbz8vitna0+O4UH8YiPYlO3gDrKeiGGyb/72POKqkkNZ
OZGMOYTFORWfsshkzDihvlmcSO3ZwBwhRh8P8VXltUEgD/7wXR5NnxUzVSDOcuq0t0h+00f3oXTb
IgYb/8Rzr55ZcopGmcGHvi5qh0vh4riN8yja8fFh0l3ha6G2+O5+XkxBCOjLyW0luF0OY6zElRX2
iNY4hmTdjRjcQ6dRAg4Kzc/HOWL8pA1lI4gx0qM1avNqHjqRqw4biFp43cNrSjmfszaIRJZgcix2
vwg3eHzD8xtYjb441+WKg1wIt7Noju/xN2Y9T8sVeQsBTericgj1YFin52QxgWo71BPjYbDQ+yJy
kdKEzy0khs/110SBplrt0dk/iSR2mVaBzpp1ECYKPdoIzZ6MTN1qpa90cPHRxy0ngjPnVzemuSmi
RHEIFiZ9nHubiGmN7LTLAnS47LmjRxWrAB6AHDgGOzkPzAcSNRqDv6AAS+xpyPpft4wnb2UQt/El
ijlxT/R2PqK1fji6qOoVaVQCFsZk7mG1hqTCpluCkkkM7krpPpotGudGseleADYe9l7iu9Fc2WbI
7GB7sasbZR6SE+hcV7q/v3lxJDVsm+/+a7O76uPrzmCA0y/BHOuCq6DELTtgJxPQPY7JQXj+VjXy
SziN+cXx0sT2jKyFJgnbfB+eSh2t2d/ISoXIxAiXz7soTDJvcmnMDWzJFVoCmMR58NC0ckjHyANI
nt3rYM5gr+3qKNFzZOsouIONpsNOYSpABI2KEUQKIyPvKvLc0xzLOxNERmbyHdcokVTvwFE2oizb
eoKhdJSsht8AXP7tP/8DtCV3y8QMf9Q1RHCTnMgatFTP4Za/DlCu1P/nGmk7tnmGfwKD/VfZYa+s
0xmBAvalg1lphhc8SyUAr7h2aEAmMQClzeNyeN0TelK4gZNptdIvLk36GFpdx0WilxwfZh0mY3cK
TJowb2SIWT+Dt313xbkf7Wdu/KTkOXoi0EJt/qcaxM49+by3cnxzwOYo89J8z8LxN+1WyyWOuoBM
fmAucoCuxKS6mZK/p1jUp+upglTFqdCVWiwCYXAx3vF+vqK8kgNDU5LflbOlGSp5S5aYXR136AeF
v9jYxkLrvLVLmS7ScVVnxFxJe9iYD0xny9mlZtbXl69f9qjN0asy4r79t5iNDRgPCt5a7t3lkHac
tdUHgejxaSUbND+gWXm6ok2yBpx3U3HhejQVsm4R3Xx6R6pDPTg8aQM+acsipgAYbu3ooSZYzQmK
H+UP2P5v9X++G4poY+8KhBBFokG/Ga4USJaaDDcDjoM8JlF37Ge4jGhvxOkY2rBIVNHg0qQuzOMN
bC87oCXuka5iBmOpfM9Alit/g8Y1fMFYzotpKYGtj59Hlfm/ebPvV59iC0V8sy8w0AnZLprs1KKE
eHDvbuu7H9Bf7ebPKpfttMghM5jzWmzNu3VOTvwbJIfYMlb6e0oi9U0DOSBem08KQJJtRsNEyFTg
R8p2Vl1qa2iKjQajO4rrOc5piDsp8+5ZZar/ZOu367ZgrzONsnAed9YZQuoBKK1RnNaAI2IzDS+q
CDuQEaqNUjXivKLZBnjeOlvA2n9CnZoC7V6ioLtiZ2u8jLS8wIHpcxwcHNZIbuKPYjDn60Rb9lrg
NiHU5YmluDdt38pupdoUKEY/vn3OH8aJ04gJB9Q91CupUHgOzY7ZbVNpjGuwRqZaVqZ6BnwStACP
LPZNRPeHGwisTunrm5Aft6YlusB8A/gWz3UWQyYDqZpK5VTkmSpsigRz5F2enBevpPaCJnxeV5ix
lsi1iQFO4T/xMTWCJh8fS3R983qpdNnpnMfKGdBc2Pm6ItpGJHtOkihH7f7+44cqI6oHZFecYS8y
ydvgEMYMxiVBAzCyIQLPTfv5ueQsjK49oKedXcbqo4qyyE6+CoczvPZicq/wffcFNTB8N4FTOpKn
QGfctjE+xlmpLW+a+Rlp3mTqVIWi9+oTpvDnF1vuWXOjaowGix+QAVaO0Ur1vOwBdlyRQF96A4td
VAm1En/kAq4C6PeIv3EvL6ZVT/VdwqMFZTFMsSKs6KZxuP84VxcPPHYd3SXs2BsuUNHDtYtuX0RC
aY05x+u5V+eEQN5oqrPA2hvDVzRZSljsjIKTniYnwSZ6IrWZXYpjhOwhjeeqkPFyy1fGJk4wtlRj
k9pShOX2i1yhY3jnqixzi7ubw3gz98AFlDbd2CIgiaPURKqi2xs+RZkfKLPc1+rxd27wjQtzuvy/
02ISCsMaU0b6U76jIHw/gZRQQdCdICSTNbhFaaj4OllHbqBcvRy5gB07sSDZqMNyZH8kJO2K1gCw
iojuKyxjjbP1HyhDHPxfWj2K3AZeplR6jo69q4qAevNagBxrfFKMduHmasv33TCmFa2X77bI5lLA
vnbVRK3ITxk711FHLynGylxr8HXPFDSWJWT7akp3qLRK2QeIXXlVUxaO2aY9KRLeME4f8RuAIkd3
2kcOZ56ecnez938NjeWW4URY4OcnOjWDBgJYhRec5sU1Xld2igJE6kSx6+Bq8va678BRMVG8MTUR
EUBvSvZRugQY4mH1js4kYMQJ11fcQVitKId1MpOpVklQi0rUEDZNK5LmTug6RtQ5mXhg4jpZg+2H
O4+SIjjOS3iEiGb6i4WJwBUHAvJodE5B2FCgRu91Hgre49fG2CRxwPRCL9bwaDB6Z7xKgILlz9lR
+4bqDIYARB5CqFSa6XEUt6Ffzbr1DESdJ9LRxwSEovH8sa72Zgu2IGzGL9u8mfGUHrm0Uy7JOxVF
SYuv+blRaJ5dnFevrj6bM+KTIbeXCgmOUZzB85O7LBpVs2QtCU8jsa860aLnqp03156l4A/uzFuV
M8k2kvZhFQzsKG74GU1bWn9KgSNJYKf4jzWj4SunypiC9vqToDolsb4CVxzK1QB1tinpgoQrewWJ
BOQIU7VOupjM1d2IVhknm9Q6vAS1VLztTFXEGYBugXdDQgSg8qDqcttkjvd9EyfPF2c+qBN7O9/J
yCyo4bLAKYkiMPYkfm/wJTLTcP8bmu8mi8aUD0WU/5NzLB+uLPxMol98czeCwemYjfD2WbIMV394
cfALUspLrOBfzqHLw6VLHamUW0BT7laAeAIM0ouqWXynIstPdNSuPMzzRONoI9KqGb81c8hkkxVm
WeCg1NXJ6OzXKX+6ut57V0B1mm2XbAhldJTQrUXx2RoAf5VWClxtHGnf+bHGTlZcz5rI+7SXlTAq
9P0iVQj9aVOPOTaDs5gioa21B99sJFm21xtP8fy0OLkTuFCb+p3OOVFHi9lE3RK6mVs2z583sdZV
AZ87LtD+wvpgmCxueN4GF7uu6aP5LpP/h9fBx4ojPn5SgcZl2q50H7B7URzcqszrhJkBX2KMrPW9
fxMxY60YXEtJmfWijIKGqNpyzLVTrUWopn4a3avrHX4chju2uym4uJKO8WFWocfDRDaFHpY4Hj8i
OGorCIN20mYqB5iFJwgzR3sZjWD6JdBs0RwZHKF28arCkVp2AlybhAJEGoDvkzdbv9WtzVzX7vRt
vGyrTUu53+yKpnT8vki2itRJuVzYhsSGiqyRqspTSiMVhOPRVRYp2SGy9p1k6Y1aalmPGgsJ0HvP
U5/lfbMLqgrTathjPAe2gpP8SjHGgJtgr1m2m7TbP2T1irE+wDH5P6p7Lu7ggKbjvhfV4iuzRYxC
A4N8kjAdqV+RrAFL9fhAvQ7eNcy0iAbCkDnb4RS5tkr+QKiq9jtOML6jdPflxxPtf4Vo8oKYqccx
4+LMzAnaDbmAriMhkZU988+li6sPJ959ZigPdMlhYsbuL1W3pmDpyb+g41B3h4+Wh0HPmh3wC9ab
ECCt9jwxCNNxLku4tUDQyaciPK+SNdPYS27dAokt2APgOhBMcAKWu1nVDgszIXIvvawWWGqRq/R5
Z7aaJr9+Q8RaOMBuYIL15kVxZ0RvYYjVGrDvelWRofnE9+YBrjPycgCil5G1UD/U6Q+p1msQm9PI
Ru++YhDKGUPcih9DhrkPB35YnCiqsje69UELElIKU/spsrxalVWur0e8N3LGQd2gFM+dCZ2cJvt/
NHPoqUH83yybK/Ak97hy4ugg8YsKuMrdaHDRcixJ/1q/FF2I4kTl8URZ8gB1Bdt3OGMPjY6SRbwZ
kL0bl/QLDCRctdyVCHzcxiy76vqAEJ/Yr62QytO/y7qpmp+Phgclm93ow7TcVnQJiz7hwYZRDlA4
ViCoUVje4yzm+V+dPxgw01D0iSQ0oAMgR4954whhFoonZKRzUGjqELWPzgzclFM5EXyf/ZHrDdtF
dnla+dxoIS2zhTUEBN5kvNJmTJy6MfRH0xuWyFevumkseoli74pADP5E83RltRq+Pr2WsLXUvPrr
0Mra3Boi/0iW5i2ZXmaXeHYWR/PUdDe+4SLH3XFbfeOv6jP7BjFwNlzJp5vO0pzefcnmK+hcanXZ
Ltr39HmgjcHqEFxhJi2tC67XTyQJirB0bm9JVMnaa3rg3osZL4eBUJjrI+XP0rY3Ef38smKvMv/c
uDKvYe/G8zYWrii3XmC3LIEzqOcMC5AUDDFjFMI9B+i3ASbCTQRe3hHp6sNb0LX7qvUJIePfwM2Z
eCKNhZsU04YghR7eCCuuxOffuCj2heUrq9n704HJSfOa57X3qYUiCumPQsiz85ISFhk//BGTiU7Z
Yo7Oe5lwxWmcKH8qgRDW4I0EDk15I87O/BnoFS36da7zwAZMioePnzt57lrh9RvuAlxnbNXhgQj2
vh33UmIHbsUl+1OUDvisBlDX0dyJcyCuazKKZn1O7hue4pexERHwUghRlmvPx31fQ5GjeqPb7GQX
NY8g4dcXSvxlneROvf1BWyCvzhFEmqRE7qUOXT82UC4+dgZT73fKFYZ9e0VjO4Id2jNuPfiATGjq
BT35KLH3Qi5HR7uqZI5QnmpmncdHRopt0O+6lBd6htL5p4dxRnwWt/2hvshvk48uGaWwOrV10tmB
1M6lDsSZzy3NGVMsCc888ix9E8vMr/IPpz3lgAtSJKj+RvWFfHDa1bVUQHo2K1jQqUGLMM1WXqCh
xEV//QySTD+OuMtoKVbShG/NeOi4dsYTKH+D7evTRDUIjgFWOXJMKMVbBGzCzzGjWmiQJe5zhPLh
1Mktn1eJ1E17Q1b+F4UkXqoCuDr5SxJSm6I4vqQkoqQ8PqpZuPCTvtY83NR11bAGVDWXXKg/ej1l
BtG2StXmR6hC+CtTLCVknCs45c/2GdKBTGQHc076c7isqKx8eEViEBX8rKT4uyDvOWLy8N3LMncM
eqtvj28vp/YBv1w6ynJ+khvsGMIcPiV/M+j3sztZsl9rIzBeQFRicazKNkMySph1g8t9cITPJDWs
z7RoZhr7KcfRI9M63PLhGvCwOXgw5okPtCyI8hxFLR0rjIrze39kPRbVSBkSmcRKRsg04g6Sz0jr
Lqw7cJwyt3l/TnnParY6fRRZvg+QV3jryQNnIRTArDeZGdpqmHVzhejUACeOhTwTkyZwaRnS8e+V
siBLtr4yThBxZxQLpm857ZBDaVkkEYwiyC27AV8Y6E0hIayqymH9cud9PayrQeBoiI7bjP9VJ1EH
cJ5up6+C6plPV3bOFj4M6hNMnT32JTp0Sg15KifDgcL1w1ZYkX2NnZ/yH8xjDMa5hgo8X85hGBYy
5NqBUutmn6iUbOd8xezPCbGa7z1OtopcMqYfqpSAKPaC61agafG32LW0LW51nK7jK5fu/qUJdgWD
RDC/8DRoXQico+ds81ZBaf+Mi6R3Za4iWL/ccs/SnWZ2sITjLt9e4aKB9Ly58NNTdvaluQTMWhxy
FsY8LUhEPHrSLIaldJlBpvEPl9UYaUC0V4nzyfsz2zmsao/2WanILW7sx12CPe9E0mzDzDWhexTV
BEi7OX60r+LuIG71TNgHHMsrFRt7lp2AJq6addDy2qLVwcgdNikAVMqFf8lVnyqHIU33gqmRS77E
NDPUUJjKJjR/gKdDN0FVEXq3ZTiJr8zlKlngCJZW9iiZRFjOMpAWs1NNKWrj02W7vcpf7sh/1r0B
G+TfbpqjuU9LjI03P5ULjUFvpzEE6rN1+/kF/s/BTRo3x69lD387OmlYTr013U6v1DdbryuhD2sB
lK2WyQMfa+Ofv+z9clln/p/quQl/5MMDpIhwbRTUA7ZzQG9DWNytum+pC3w1vj63wILobt/d0Yg8
O5xmPCGpG7e4BH7ZiArsxzvK2jy/QBa6ZXwo1xR3Wz8Kl3ciQ7H6fdDMCxR3dhBM3khNdRXJVjLf
TbLBCkpDrt5kS9eV6yWeruN+Z9pBUKB/HzdEzN/L3dHe08M6SQhR2UGszDd8NJbopQWEpj+mIuy+
3RTvF8al2cFYTjf7bhhfPujmOXZJD9MYvxm8r3hsnV+7ZujdfSHOgiNgZjydIRS6oOnwHAqdYd4X
Vv6ttMsRNeSVia2Bdf89mpVETHS87o1GwKSnceoXwEXHOkqor3vvkf0a5f0jaa/eW+eiHXJGjYk4
BX4uU8x5X9rqzFeiCMH3GS45S98wJ5HpShFNwNExdCgIB1L7vyMA4SrO/IiRAOcjfL7vw0BQklJN
nF/eKiY15ZXsivbwnFQ2KtuIyyojStSOwI2CdXWOHlfD793ntTNvwGlwBnvqBO8BmcJzYQa0aiH8
sVHDPZdsJxwsEk43eruebWSnLyPgVGuOCI5OdmrY2EIQjG7DzDcIbnSOzFikHY4hWLyLKJkEh4Z7
JIKPb3QF7PBwzhfGNl7yDiyXf0R7Ie3aWIURimT7p43PZKgsrNWsZOdYDz/s3Kn2OwLRxZ+WJ6nK
gMIg4hd2FnPi2LAH8IrnmaqBgNbrM++8ACIkC+OKLGiasf3SLXUenATTygI1JVfWGfloprInp/CF
ktlOnIIDOsEAey6H9HS6s/0RoHv4i7V0Ww7u3DCchI1uoIy9Hz35fTP8TdEBLqAZi8QnfRuEVB9m
oLPGW9KkFCd3X407wpN3YeUc/CsUyFxBfVYW1g+RnD1jZJhiCcWtrf8iBUWD6YP+dU/1dmd0V2xt
YoCyLA3PNT4NLt69J2japykFN4ThmhKspUtlDsQChFDibKW3HJWpHrkYLvkif9wji8Ophd9yTSi1
sMFB5CSr52dFSmIJ/8FTxeFNzhPHgUuOHvsjvSftu1goA75mCply+FhRzsa+6bUnnpGhtCNNfw7e
tT2LpklHjjVqcxseOEnWxJxgtEfXZRMM2KgdbwkslVyWhYEj8X2GRUV7288Q5zwQA0wCvmGqNhzn
gm7aFOzVMBU50scxXL/MyMJYOLiE9haBCR/9ha9GHgz1DajBOkqs304qUQ8hQZvqse+HsDQMu7oS
zd+O5Vj9pDuezEqXIw3QHPQtbIZi6ePCFKSTBxxLXnvK6zUcjEG1Mel8BjvzbsQ9+EZNqdcsNyuK
ufEVflmEkDDwkyUt33sXK0KEkMv3a1jAT03mXpvQakkGkQmWCeVvQZKlcGhdvnfrOQaT1SEPNirc
iWDR9SJCFYcnpaOvVw3SQmTcD2EUUiTAX0cVzMl8N68zLk5y9MvTnGFBZvOpg95JrHi+taJVG6K8
idb7Z7roEjveaQPnmA2V1CFFCz2zjIxt3IpYw3HwjhlMXsJz0vMxDItpGFMZCuwNsUPnc0zOo00N
wAvJxEDgWK7gb9o+j4Kpf1ziKQKCVEUSQp5JnAr38zUJnnmCENuwwVojobvTyw88XLG7HjsQks2C
iiujoBTEg18jgOs8WqpAQML1jhuVZsI8m3vE/HaoA3p3/D8t+K1sGKtOndixFjur80Q7oyEJoLgH
FUZnuxV4FpF065q3x8TuPDVpzhFOPmmGcrnLH5fsQbI6QMUf4H0kWW2K3boHl2kD9bm5nGKg9kNv
JuV0gz+t7LpyJZzdDQiNaPqbg68Y0XNoRPPj35CwnfU2FR82e1XZb01k8iioT/D9BIiE8ucHTjaM
TjvdC5WwzwNFWmMuY7VnAfnNEGLgreDvDj5RjermtTFR89XWWFWi5n6nV2b9s/oysmQGK9v3nefD
YhTdMrPcAIbzuzQeKSuB7pHjTReO6YdqZkcsmengwcosQu6LJbCbJCDjekplFrzVWw1/JN3CMECs
sHu/76WQrrLc6ixLHJ3f/dnt19E8Qwe9sKynbFN5Yo+a7mG2x+1YEeFU2xno6DPytDqKeUktTjqX
e5cATY1jNqeSAjDprzrAEQAG/CrHuEKQ2ymvoqEnel5153a5//w2BgF4OtYVuTyhIDn5+mrV9dwb
Fe/MIrqs/VJzHLf6BBKzvZZPTJ9CsH/9AX+Li4HhC9XCbkpR/OAmvF4oj2bbc/D1LzSbsMToC4m2
uP2tZtfUBDO/IBV6WyqPW2WW2d9g81pWjc5zFJ92dLaDBhFn+2kBNf20BDky1LJedjDdgAkEcRK1
sLJQ/VbwY8frmlcb2Uzh/n8kMwMFQ74cX5ab/W1aI6t4Qo8/up6KR8h8MUSg1Y6ZrK9MMxOibA2G
PL3dOMh+femQ6wu8tD1qdD8RqLRcb3bler5MGESKx+/4ha6hAHlA5ovKAvpGK/PDjtG+p4dY8hW4
npPspY0H4/Ji5G3tzW0M906vYkrKOWebxgJtK88ea2GwTPX73P+wESrXqvUMQJ6hsx4mR+69M8Ao
w1Gbo0IqXmgd3ugUrUUh3gzmxFheMMOCUJjsdhJRORbgARa3/LOgtKx66/hD4/FIvsGh6H6EAelC
RNz7aGGLQpJ14EM8J75XIz9VIiH+Y4KxfKdU6gr12lu4vWBt330ujhIh9sMkwAPklL9rKsd5FveX
6EJV/WAPQenMJZXDb1sNl6NPNz04cBtUJorXdGn8d5pwdb+6HbAnHBiWO5axVSsIP4OC4jRzr+38
RADN66dT7HbEppiqUZkj7qTBwMy6GuouQWieDWbJBj1QVsLgWxBt5PvJ/kxgur+XWekutCUTlHUG
s6gpXsqd6nz3TXhBCVJjDTz6ixBs3LwmxxOOZ48hUxQz4Ux6wQ4Gy3V0rk3NUjgw5BVm7/IT5Do8
YuPMup4puCG0dRMYztLFBGFpYPVA88vuzjY8+eS+/7nVceaPSg6j5nM6ngHauWp8Z5GDTVJA0iqh
7XTPYDCl5hoN9L41z/kROEDBZW8I2+G2/HZdf9kvr7HpN2qv6f5ZIRfBSp7JxncLeemGoSMfT/Ay
yU/ZllqewDYKxAa2gZdrs8FjtIie9voL6IjNI3MiNlPxEzwQL6cStQmi+WV2DTQ8CnOoghfvKq3a
slvJIbmulym26R9w0KmGbNPUUiK32E42zh53UGFadrAeBs0VCdZa8Vmy8yg86orFfjCBI+lRiUvH
OYd4+w/aergkFJZ8vFCk1sX7m8Q6jJWOA/EfD79GENWqVI60eH9kFGkITlULbxFvCiIKXOYU2d87
qe3YHZYH6Kyscztpf9/If4EwFDEJAzKW/XJ7YwKkTaGpcA10oJ0Zz3nmttzJLdYWT8j832zncLQy
VjUlhGAG15gdjYXCcVxSoGhBRhpkBRnBt9hdXnuVKPqQ6rgFvE/ieBmGQSGAE+0Q9X2bXxJk4uPR
o9UHKMT7b3TT015ET9ghXkp8UF8qMK96Av/XQRBXFICEPxMM2AlGjafw+pHxEC8Pytj3N8eCNho0
6W5N8xeebuqo+JXkEGqpFLMZ0jK9PSYnsFiD6pfiGJLXFrVbRPLLCTfjqAeOaj7H1tj5hMOC9TUn
po4im9zgrrP63pYNqRuw1Ts6d74XxUIQNxmjZFWYq+0tbcBMhrNm2U7rvi4nL8GU7qll5CiR7oDj
81R3LsAczgGn/3ETocJuUwjgS8Z4UAhl/oGdYcr4QFPV9Q0xs/Nd9/Jx9xPuadej01sFJ1JIP+19
3X9+xVruV/Ue2Hk074c9MYkyMH5i94tv0owm+DsuOfQQLnenCDRnrDEydLpYZgV7YFb6wjQ7OxiX
lge/Ioq5KAmSCHAJkOp3YqWqe7T3A6dvw8KMoi5RQRxQXcBSjusKNfaWDo+Ita8Tk10E769HM2cK
SAUQJBcpbR3+DIUfa/Qq2OyFOpGsah1cOXLedDyHQ9YCMhrepG6D0LNWaYLhKRA7kdLxwk7YxwzJ
D7Yw54gZSOu1lBbLWcrOY+rTjwR4Nie5loMY7FgXnBRybAAb2zohw9xzCUWySlxXcsjdXgBoMLaG
119UqNQ+r5+CL05U+S3DuHNaS2DcbY/NiEOdCnQOYFQUMV8KBAle8/KU0vCWpNLkk2/Q5f4osHXo
0IaXGMgl6GGv+lFSxhdjEQP9bUbU8oAh9P3Iwf0o+5/X5f03zAlZuj1U1O805iEtpd1Om3pt9xej
rbVHFAegluJF/Yl4tWTQwSfSsBgf4ySTjrSnd8BoOyrGJQr+CaYVnbru25j+MyzZ0FbsaAS+EyEK
5hciRwlcdjvpEwZ5NPkjJGfGSurUZ2beYP0Jj0/T6iHTGRdM6bjUdb4IndvmkGYU6HhesVXiZ6K8
Y844yaiZBEjl8GxFzx73N1QuZ5tFxwd3sp4OF/lhORqGrQ/4xlWg5SHCt56FwfjNMPJ2tTFi5D5Q
jK4U7JLQNJ0skkD3Lu1gG5gw3hr+zWygCfWFLVWEtg9WbJWcM5qFRxKqpHLqN/xrSvE1fjw9Fo08
L8FgrQ30mIHk8/m4JpDahFk2NijyzRBt+f1GKfuafWhAnXYjWwFlyv68UrhNgCe4w2Ioa7CFekMp
WiQ/aoT0S2Dqy1+ZKU7yI/yOU4QNxwB0gGy9Ch0FNVUDcuhSs1pePuBQES6SjUp5CWQtZZPH/Xoo
Kb1O7k7RCFDm6Qg7o/38BOkpAqwJh7o8LUQCXO5bequkUXzQLnCBphwW+LmvRaK87YM75zXPh4I5
15coxp5rGjSuJrJssmDz8jE++bBpXQx1L2WzplNmAwcebTspK/UN6P21Z/L0Wd66ZKSjcbutrrXs
/XBPLwd2I5oHrMwYoq7UN4lNPgNjhcWLPWN0zNgRgJL6LsLk5QH67xihkAIe1+7Kc+BkTA33pxNQ
Okrp/h6WiADeigPqCG8BLnW0j7s6oa5s4z+KJN0HVi2ZfMslW6cItgjXX03w+zQBaI/0eUZSjvYn
cw12L+2xVWMue0M2FQMEvViJm8A1P7KMEpK0rVWuO8eexIXA8Ut5Gp77aGCaKQqGnzxThVLCpNgU
QaFoiNQDIimyOCIQTNSCNXouAlNqtciK2OagRVmJlnrU8PzJx3K+u2qmt9I/JOrhM1Kur/IONR6i
hSm/dIEtMXcnX/IA1d/76Vv0EEWMwxk15fZfPQMtmB9FD99QaQtS7KzI0pFgeCWtKr5KNMfYcpds
6suNpz6+eDdejYds+cKHyt5DSYrJLS1Tfuiy8K7AJqRsH1//8JgKJBvRN28abGno4pNLMQHUuyMW
pLKaK8ho6gQahHR288LVZvVqQX0p0F2s7gMYlGZrFQlH4XhgyzLFr4aXvA3wATXk+EOwUyHB/0fz
CQt2GTH93Ih2fIS3foRFKZP6RzJavnXlUWPaLBV2MAHSueoSLPr1ZfZtH81ZaAV6Q7urnloVQWZm
5ar04BwQieGuvQ3PFuStmSKHPTzHpSUFPKHMU21VDoJJOoJSG4e+K4jowU8fFqeu0NSG2k+/YPsX
F63jTWIz4hQxcCvks8aPBTYxQpF0SJLe0teDvdQiBlxuRF3eXtDAd50IXEMe7N+XZl61eQhq92IW
1AFKkzdK/kfSiy955kjlsstIAIbyuvwKM3YAxkGhQ9oVhlQw1BWPqLcwt45If3vue3e6YZxaMMjG
KT4WUxtLvUk0IzyQNHtZpimjKCl65ojFdnU9GMLTvraYWG6TFKDbWMc1pV5o1CabNSWG5ycaRR/W
xxVfAcEEa8I9917G8oiCFpo0WYEBcWdqU0/sj5PoOp39bbmo0vi1MlKBUvotYqCLgmT8nl/OBQeQ
fmMwB1+6eO6Ps2cC1dT2S4JfvbizhjT7QCe4MsXILjJb8BR1ssZejgsddHtzmbZs2cO3E+l00bgi
eg4Ur/Zz5/ftMUsR3mwoKMMFAhE0o4AdOV+CBSBOwF8YDHF4HhB0P0G0JWTQengT9y2/91kx4gHD
31kCoYth+jLMxMoXiBMmMilnuV73jruipQaWkn8rgDWxQTY0KriQGYWWea0F45MxRZa6GpCqOG/B
iAglj9FPUtZetzYB8SJGSTOSSkLjbFBSOdc9YpjJtdzkSAhktr1AhLCs35JAK4naOJ8sWr6mOHDY
0T/gqlsX2dWxFyEtgkLzc03GThbbTYosgPeOk4xWtdCPXkjsCsRUe/KPI6GUwEPWScspBw77Vmjq
OOmZK820weYWJWnN2jRUkaZS8spjebeCCvSr06KxaBRuuyJNEk2Ka/GJoglYYG4SPnljXzNJSTi0
LD74XylEvlHZz1dH7oo9fRHVPPeVkUoI9GdwPDPzKx0Vw0DMU2cdP63oUrR6jfpgpv0wz3xbSNsK
2OF/BbIOhxfCZVPJJ3pQiWQ8TEyxEA17MeE2z6YdB6aPhEhp3MvzR6hkuw1/6d/cVvA/rD6YvRz5
rRHkjtwybbkGm+A5RvHSgllLJftseziFr0bt4ekrCoAE70f2tHnW78BeI/b4qrAHqquiqSO8r2Sn
qQYPhtGGFGa8fEfdgN+/Lyec33yAO2J0f7kSJtGOZfGdeQWzLIUkoiWOzY0gZ4vNrzRom+G7KJye
iOBpydkdGUkr+m6HsC0emPTpJHu5YVTvSzx3Y6Hxs8VffAXYdAkw2+ZEO69bRmzzfJph375kp3hZ
eGIkCqBopo3rG4wss7zWBJ25f6hQYuGdsEOaMiVLNDzmOhTbbgRgdWypevJqmIsccZ5KFBwETYpd
nwo4fv9dd86tBX8GDa9Ds9/n0gYLDfGaJLKGAoInNtDXEkvUJmdqoYq2V5dx4ruRuXXZYXUxrsNo
UTTGfifOK7XSMAyOIb4uzxj+eoindH+398NmU8yjlonRPZ6ZhqdZ+6tpzy9DqQsUwwgw512oUTg4
3j4+53O0nmdvVMOG6jWZpitEfO1t/khgHlzt4d357q6Q/FVue+VtnEDZrCqhcpi4/jkQukK8PUSO
AIZKTKsaALea6CPrQfnjycie2sU25dB+WqnviFTGjzb9rugRFq8VHUfgPlVWhGYgo+fYe/OJZY8Q
LT0R1v36ozczY3Be361uTr7WL9o69CEWv70UhPyFTDh+enMh2Vybm1ZiKnHKOvgp7rw16zLHXJlH
+zx2xw9LmLJgmATVA/lHYTQHZuxwwhKoNLwoMcDdcBW8Un2wxAe7VukqM4/2NlmLkKpYyxCiKODr
5VQXfaYEloV4+uiJC/CiL4Af4Pmay1LzJVDRrCcLwq9t1g0TmKj7bIucWRt5/m+R7vzyWOzM94TA
BIFUbUiC8Ss1HTljN+rpfHfKp+y1f8y4UTMlBs6B9zf6/9QFfsofpUdY/P8T3zbD32OmFBvh27Xl
gBsvtKoG2h/5QjFbqCgiNxVFaJf1m8ztGyr1e9r29a/ugvoGVXBS1CCLitLVvLy4lUyO5REt7K5M
mf6+8h+NgM4/+Knsw9cc15n2fUOy7LDuMKoEl8QPwC5Dd/NE3nl9UvPnEE4c0FxLVa0PooeJsAu2
zh2+OziVnvOG1j2pf7fPTUNDfcMcqVo3T7bHd4gPuTCPOeFmIWZPWZo+5jK4JT3QBpydZX81CN9x
iknc3U5bwo2NZ19v6hgahRQGHy6b3lfftnaMYd5g7OxMCLyYMVgEM6mzCITLWHLXMVCKbUu2SgVZ
dF5l2t837yRJWC5svYRWYOwMrrf9SjuIplgeGZ1bmqRAbePYpjohnh/j0gnf5U0eAJT2nEymAww+
c5xOCexOca0RTpsp1W2Ed5EZlHReAlD5wz/DPw4/lOy4VafqPGAXv8O+7Wc8Ht9qByvFfmuZkn/6
7E2+pztFplaqtV9PHEGhkU8MH1z0PRgtFWXLZWXcsFOLbgOdjT6fLodVQX6xhe7lLB+cVtrl7mSM
jbpkslhmyRNnKlR7xNVd2oU3FW1rwwOMNEtDPfLDUSags3P7Mt4gThhgqLwkCqxKn0dNbo6WaDFb
QKirpOpaEbyT9mLzfQVKPbCjP40qPahPhZinC07JYWlE4mycDaZv3LkPdkFye+QkgaaQXzQHCXmH
wrAveYsy5C92yVY4faAbg438+UzwJ3IFS6hzAh2+IWfF+oHjhjxZ+5irlljK4CW83eKG3Emb2YPM
R9VsLaDP3a5805fR8TP4maLnCG5DVY5B4HvHXab2pliNP2qA0zVSSsKJZpqDYYhYmGoKUATahHQp
v5tjcoXS2rDXh3ZRVfHWgPPYqzl/F64P5EFzgjQ+dmtDj9QuuvLaYtWPiBKbmrwCbmG9nYEIlEZu
/oqCOUsr7z065fsdnbGvRAirYranpyeaNFKuRfo6qIQrrqqJgx8Ci/qgNYHcZnqDmyP6Ve3iqKnx
EAYiCwTcfsmocdEZKBQfx+Q1CO6Cfg8CJdgU9ZTFgN3bpzJ72jSB2aBnc46xGlaLglGUW0eZ6dlB
O5aw0nVrKICPQNNP/WlPo4ubY9DQMF8JaNehOedHutcFAgGBVZEPk1n7fbg65TEKb661z+xt2kuF
pJKSAjlKV8lB0YZk/UQ/q6Z/WtkIuLgASd0uxipkPSbYnehqu2g/o/XwzuHx+qCu+XD5yOpjwb02
yFHPlraW1f8ejG9HSMAQSOJX0MX8aBFhC085cNr/FtkLh8xjTrG4aPVL3/VvmX93Yl+laviwnrr7
LpiDq0sm9znV/eVCIRubJegeHBGmuqfyo+BXdRgmiLs1rF/9Xs1JW3bF404Dj82hcfQstr45fDwM
IbwNa2FQEZF7LvVc5F9OPikXLyyuQVAG0CXO5im1AR3jM8axjx3MxiOp5FQ1n8TI2lpwbyFh3PrB
y/HRBHSgwot6cdQsP4UiC7dBP1RLV/E7U7LnGiozUNasp9zwb6L/cfdj7QZ8giiFesmLBIckuEz2
W+vQnn7A6o3kMOH25K/10xw4C8gLFFE8fzcMsRJpByYa/Z/bU1QGsmZGGTdNvhu5aADTUfL3Nh5i
rfQsQXM/GPHN69iEpIWXRZ72vc2QUsxrtIup9SYVp+vcdkg+g3h3XE+MfXNX3OkjHf4hpbBR2Dqn
33mYrvKnmOYaMPtsFK1428aOD8lp09u5M9oUImfQUJoErEhEoyuODtbkrawChPRu+jwvX4pWyMae
AiqgnZ2GrsLsLroO1EgZhISAIVWoRBSQaNQ1iHJ2Uz+59UFiJaEp9hpwAHuMqQSnMUDmIf3DPYTS
jvW99cbsKYYhBaCBOMIVJe4XWWQgklKPXpwPQMyplCaCG+NOqHThcv/84fgYWBX1klQ4lUMVfPR6
4WWVvchzLAgTQrWs0+6i4eyuIWAQFIURYWXi598CqxcvJx8mGxoIbDstqZXmdZMwN3G9Hcrxu2vu
Oltq6Pke9R36CmqDvt4yy/pYvkFH1/91prdJreW2hKlUzCKVkJTenqR93J6MhRpd4u3YzvQ/U8uU
goDn1Pn0ydUTCw25zw3o9Z9udehBq2Hsj1QRW2KJySPpA8k6rKXLr4oY282l9LJTGdkLYPyEQySD
uB+WcpjRLZeDYcJBNv1Xh9Nruer632v/MDJL/Q+Zu8MVApuBH//rcHyX99RdvRmlGl9RhemBZfnN
6nOHY/um51NYzOJWHHRzsaxVwJbmWCfQGFO3KA6A1xnc/LX/XTp2V1cthSAgQX3eEjj1DzJHRjza
MWDsfhAsegjVomSMp0tYs8xZLW1BPnP0a11FBsbI6nGw6Vo47sTuvalhd1Ybe3u6UPJefv/sRG0w
RctSvlQOwgCpskDgSyH2g+4BPmV4pIvCJ5/4tnUq6HoTamzjzBMHFVb57/jX8PEHh3Tb+ki26J7g
xJ+67KO9CijaejxVNP/ZA+Ug+EJK8B8CO9SP1b/rj4SFfAaDbJ8I8QrJxg3EH+GWGHKC/Abd7GEM
mh5G5j8bHZ2NaqwfBSxO6tjUt2xzElYwmBZjRwLUNZH6eHaIq+rT76JVQ6PC6iOU5+ydVnkBVV3+
PAG0yc5gNDfE1iah8FuvAhfuA2OnarPrLky8CTPfxMf6t02Hj874N3M/OtjFjWvn+O+eZsOSHxx9
/2Lw3/m6uNIsqCfIbpz9wkdqMx5yHnuBN8fELWJRUj7u40u5LxFyW0wCKWifZuUL/V2FO1vjrngj
hNuak3qSw6XeMhSfuvX4odvaorvL+9TcvOm2lFWAR1Xaej1M9P5s/jpExkoUlbNW+kC+TcJK9SrV
AhIQgDyHfcAq2MK+pZ2reGDxbHggBN0RtFQt/q8lCaCIQqC4C8f8HqLZpaaA7lNjIYxyv7bs7yyK
WpQVuSym+YCAISM2jVXV1C/Y0dL09NGj71q6lH8wt0e81M4MJ5GljyqL6INPbK6R1BXIxh4KRJJX
BUPoBcz6HOGfEysWuXZye3JLG6o7gx+9M8YR+vMuS28YHs+DnEOh5ntEt7L6wPghmTnUZt3qDxku
U7fEu6QJeO0dWSsERhO31/OROw73cnJuKZdDUVR5Pw9VItNZ+Sa4us4CmY7/FYDj5PjoK7SbAnPn
zpfJQXxDA5yhvFzXzZr8XLNEIV5pp0qtm3q7OyVoRweIzuDonA5ukiNqKsm8GHXQdv0zQ1A5GwN1
0H+ZcGUfp3xnBUiNzsXj0Dbv6xUj0czqNBjG0XLuXGMalXvwuGvIk0WTjlQSf4Y1mqdjezkIN64C
Y4R7W1y1w38fdHu/zn4iNb+Yw+AnZ3LQTit4+ncEtkD5Ak8aaXzak4hek9GaXloXhR9MCGdd306K
kYHgfDA7y6fXZ69Hiby0ZMharnXtBzoW+OAwgM4N283+0EODKJHAviXNxJ7AxwO+sCCD9ynadSqc
3B7IJhzWzfAcZBMMx8KZeUY6E4jo8E74vIjT79NKkrfBmmhZQ4VyPZSGjeXkJnJavqrGRVgfSpQl
tApyoEhxkIfGPbxO3zpIKUfMy9SwTVcPvzFniNKOR8KY3OdlpuIsSvvbuPVPZptkZhrTgbWS3MFi
iRibyEzg3l7VqMttcRlmQ8qOdY17/YGaPYkNGjM5SuF1rPQKat7jnxz7dB2oseeF1yLnegXiU7HC
u37L6klQnlTUXLeXbwNBUz6JGtC8UVlj0vLvY3XYKBHMLaFSXhGagNrOfUrv4UmPaiwE8syuc6AW
TQOGsgB8tFadSNurrNuxFfdtcpItGdhHqE1uEU53DOU40/RHi3zbmxcMigqYqWKn9gsmqA/bfbRW
BKb5eROOjpN9CcuQPgDh6vSspZXKZAFstzbuyVe3ZKMZyTxZcoRo2Z8PelSb0/6f8UQ5wwnpCvJv
8/OriR1+2wqQtv8LbKuEXNgH0S2ylLxCtYI7jHoTP24nTcOpJrRauIsgKK6AgwuKsKYTFkovrrcZ
8YCjw9cG6TwToSail2+kl8dfpJMqksly6upkQgAOdwueSjfJVOZlvgF4LK/jsU8MdTteIUG73qV2
MIAXiYBvykmv/3wjOXgNvCNGpmu5vyLN2WwgXF18Y+BcNqkz+eDfWIeWiHOew0WmBGP4A5/AGalG
r3oLB/7XFpec/9Mzglc7vHYlvaXOl2w4IeOwEp6QyZ8KX0g0lIZ8MKn5yU+LeuuqUdtswfvdaqvo
a2yW6+xpNwa8nJWvjRtIhsUNCQfRwGmZZAaW9Y8tdSmSdaFBgdFSJ2ggpFOSZSCGPV0IJSzJggZC
qS5L3JqBL+0V0sq9ktO8I9MWTdlU9SWPJZUud3xzXdQLaWFKjdKhX/W0tObtxMt+/dcXEANMVMd1
TQnDvg890Nurr0j8RLkTKX/pfebVUnQn7uWoCEuu3YTyQL5eeyW2g2LyovXULqCKTNsERriBbbTb
+6FvLMnXR6jiblr1WwemQXJWmopmNaT48LvH5KGirgR/gNpg3Ph0nqlU92styCuqUtCFonjIj5Q5
xLMN7GtBKOYOcBZDmb7OgVywvDxxJoxfgFtbJBVvOGumTm7y3DgBd7clFvUDgMlfjbrxaOrTm3Ia
HJm3uhG9BKWyusQmSjOvMIt9cugdP20asS8WQUBEY2QhhDiE28elJfA1UjZgCj5pH70wFY7d2Oo4
oHk3nhAugfVCFw264DgXAGy5DeX39QpUBbst6zaZqDzKwec0TiytAyiFtEX9n1VtHaiolOFboal8
cF72rX9Af5i/09f589Doan89/188KbIsXQQyy9XhF747im2ktTP+JeeQorD9Y4p/qFzig4PhmXu9
QWZyuhDtUl7kHKWY+y9VOeLOd08Tqoi6IZLMozl25oKJnnW0pXAVPOhVIH8EEna6ZDedcA3xJDA5
DsxWJ0P2Q/JGsIoGK8eL3eXOD/Kogc2un0PyAl1T1dCPqBQgx6adG0SLzsd6NIM+dw1f69E0XVeQ
b6r6FRi3QWcRYT6HcLGsAJvxvovY33TvvLvj7bImIVYDuIsCAQVv2r9cEWWFCVr70AS2yVtP43z9
GxD11LTB+cig3tBW70ANUoMRfEZaBhlr6OzTEryB2frlHVgfoIvkByyexWLqUC+Glv6+C/JZEEe5
Yx1/SxcfDvZnkRGkDA5b3smPLMn6kHo508ak2HFN73+W9Lv6A6qsMB0Y0RbMNOJYLBut7jtH9/QJ
BHFRbmVJNwsEnYaVuqdASb9EHWsdEwfO4tDkGBTK3U8ibqzrb6l5YHiZxbmiDEMqqv3oGwgp4MCc
TgMDs8Xhaf+ZmFwaxBmBQybpzcm2S+Hum/hQJ1kvA9+fmZB3RpmMhmOXp5nLJg64T2MwhPjZQOnO
SswWXNFiXogla/bXe9b9r5BH70dP2UVo0DPFJw8izm8aEGqmMdQSCjbL21lULexNY1pFpqWapcvM
6K+6m/uE7uxkxqduFiqKc/to1uPO1fYdby7PONu4cqMXUxdkb4vW+/J5HxJnAzBMt/ak4KKlERn/
Px91WIUUGy3jnNIw7/oe3oY/Ia2m9siZivIPE0lPgKQPPIZigFbsTVW/vQTfQ5btqj1uYzEHE+Ga
VvkfDzeviK43Z3T+ty1XznZz829PzDTq/ytSOnm4Hgi829aUR5CaIThcUFR0RumWxPsFOjfJvGs5
IJQx1I6C2Kht1EJWecfikxYqUaUTD0TymfP2YOThhe9O/CtViAm/fZNVW/VpVwgsXbI+//cokIwD
xcRMqJdxrlXOefkbO9OZ9q3lsZt0tSJwb/33w4MDQ0qksAMd8InxVF+D82G8rM8fVclYTGvcMgF1
jRGnVjppev52Gh20NX90aLNCrYvmCBXC/sAo/GdCmhLzSDemImj3wBKtdWmmtoUjd61Y/+/mVIZU
2NtPSruMBHJd5n6Q0hFctFcPf+oE+Uva6ckJCafN/jSK1kE+ntNaoK4VkDlYX+IB800Way0v1cdK
S1l04qbGseOcTOD4vuGgKB9253thvmA8XWWd52KeZf7Jf+bO2pAZAqtzEg4pLVeHGazatKoeH0Nm
sYGXBUWNGDiOnsp7tcBfuTcZDS5e8kOsxD0mtpfVP70PTJNiuwW2MVb43zf40VGDmUfi2y+fYkOJ
b/dJdfWNrBF9cVdJHxwmD4420msTw5Vsot06DY0ixABZEjWUsRK2wyk6tIcCfe2Iws/Kt2bJqx+s
CYtojjR3qcWok3UjrbgmoUU1f0MYp5evcLWNrhHkkznuoWd+nYK45i9IVOb4ITFGg91psHA7aPDD
ICAQaa12I0PnPmkg7ZTMM0rQehjBeQ3mbj/Ua3k0/CB/YyjEqpdED34CumXZF0Uwwdp6FLPSWEOk
xam0MBnI93ptwh33TcvbEqaw8uOT1pJy9pMt5ihIcgAzKyTz7FWMODRY7ldGlbkUAjPaPpBk69HZ
rDDYmzHWlivRklPkhx7UgJ3wNlV4dt8zfq0egtzpQZ8Nh9eaVh3ZlIWrPgfj+NoHh9RmUOLXZTWV
DcqroIuBhXTsSQAXZjlg7okOJgr0Qq440iQ9QDr5t/VQwICh++gdEm4QdOepovvUGbCeHRbM7WOL
LM7ESGHdEiEsWgVRnhgryQhSRJI4vHTU7MQ983EFTK6mvK7r3f4umQyNCH081DRo+vOFRbWOmQoc
PQfTJ2+ymx8JCWjGsHtiHcLTmFSNjDsdoPXD1NDWbs6s6QUV/C4gpUrx6YQI9DwdT51mJikyKTMx
64vG4YJrNQUhIUz34wBAknR0aYSD43OGGCmqBdXzipRIZfg3rSpFdZ0XeanGh90PAn9fkRxl5JIi
EXA32fOn554OSvsclgzf5NG1coPs0k8eJIJxXOTtjfwvjjDPSpoH63PPGfWuhalANIHJXrVNaz71
K+eVxl1ho1druBYlHKVztGy6W0l8xpQuVQ3MjIZt4p2vH5fdi3D0I1BuYF+vDRtV5gFA/fhrWKXm
CA8witXr14Y9BTEKZFYqGzFkURJs5+2teyE158I0SvPDWVt5fQMhz36MspEU1Z+W3wJzAOGCEXv0
m/sOz8r5goFRbM45nUnTmGpGPiBSMrfH3GEuq3AdVg/ZxT2qoJBc4t0yXGr5koXNug8iu9lg4Ifv
XWKGvQnyYvZPm9pCJC5rEMLKU5MxLtbGOAywapkdchX8AIVS0EL4YVkRYhBDFjuDxZLh+nJlV5kr
/lpGtmNSXi6UvayZ+twY9yTPn6jWBVt6Ckg4d7iIVcrRtJyZaHsuspGj3e4Q9jMVK/wBbGrKFHQC
itF8wXJA5GYGUKBF5NnTvxJKiiiKZN1wdd3LzjRdliAYcllNg887Dn3UepyaNwc5HkVFwKU1u86V
z0FICkmkA1QBNbQta+Sc3NTpqNsUr/wdWjBZx4uB3TiiR7PhCz+0LuXH0kOfLXwSWfe11SVYfLaq
PGcFAmJnO+4ofTJsx4+SCj3hi/jgdx6RjP7J9cJtt1NQlShEqPwWVUuYPPTCjuJLbnIeuYkhozzB
o9BlyyOfqSdTObti/9kCtuOfetMbHgMI39TnDrnIyJ4AiKQjXGE8F6M+qn+oKIck3l95fhXLks2G
RnIHLSQCwut/vxkB/6TcDR0IqhaBM7zLDHPUY/WYSBupxyjhqnP92QJk1ZdFFwu39nHpOC2rz2dl
VX7BovmOH5alGDSUtnHPqohBpKw0bbHaqjmX0FIaFrWyorklLsTUEu82cve2DIAO+xpwPwfkH97R
1kwhsnYNG1RuRYNoZboFuPEdUzQmHfBPJpIVuBUT+9TWA4tiEbA1KZRpRtGfsR58rJJPisjE3iCy
5UalvVgFu467WP/nHYf0RkKLo9agDjDpaisxc3uOnlVmh8vRBmQ7kOmN92M8eVYGyaFrGeWiUweA
Faeoku1AGmFWLUZ2zet6us186MvyKq4vBUlN1Djeox78EvCAkeby+FsSaZA4G4/TGc3PSm1oFTht
uwtDZmUpmTEPx8h3nz+iwx3i8erdw+JuHxXTUewtRSyn4Za5cjwgbvte1Egdc8IfrA8sg3zjYJoc
jSCq3S3XD1SbmP7TdMMTorCpTVbt8UaLuqsN+hWEXaQpJZlDx+v1Ptols4osdZXL3JZ4Bp0VysFI
dgUNuroLZ4x16DPy7tzI3gtzneplvh+U+HNVPXNvULeee0vlKk+BlGiHH5tqN3LKTc8jK+vU6HQh
lxB1DP8Zx7cHpQ3KzSoJ4y84nbSDEp56WU5DIvICAgBfwNJuBdhfNuzehfAK13/yPEbhtestspaj
XgnU/Zlh1uQ1b++2+h66eKcohBeL361rFkl2LL1VJixIi0Jbjvl3AzgIWTavnH1Q6ph1xiiMjB/c
1oExi5eOWlpgAGgwGF93iIGiSynZ9w0kuU8p6OWmlBNpwBZdn0RY95V4LD0TOQ5z6ZA6wvUYWJK4
X0mdoyPZWI+df5+nIw5I8ui8iPI3IsonUZCbi3gxsIIRfIcI9GhKhvobjnI6n9sw4tUixP6C2Ics
tb8e9XEeFtvPx7UfGfsl9RFidD5nvNn9EG8A76jHkn4U5NRDKgDYLIb0ddPdlY6iBv7nUYJw4W4H
fh2xMuNTNyWkMu1ogH4Pzp+64KbwG1m7eubhhoZ27Z+UWam6fR+utiS0Srx6ttyv7fW9oHputybl
td0l4ZeWfNKAMFSwNLNepKjq0C1p/alIyiAgyU7tbi49xigQl+vT77FnhhedWPcV/8U02TCCF+Vl
MOwlTCFTITPmqEfvLxxMKui++pWFbvX+kNZdIMXKkssgYxz59BjcmtVEhxzS8YVeK9sgGPc5F6DM
HloVD3JX+zViYRR6iFeycpenYz9QfZnhq7hdROaR5ir/SkpndZ5Kdlp8wvWUJxxgOqgh9VN1a96K
v/yV3Dhy8BSy5bMw2IzN4nWziHZ+P2GtWn/hb+LOzR7wWy2pmU7eEPrF/4KNlVVFkERyoiKUDGoR
33DPGqZF4i53WUlsHBJHqibwXC1Tnck0kpnOftzo9wyOzXLDF1cGU38m7ab7MCgSMssN1HWcO3Gr
TYDmekadAzMyHDd91imQAdK6Vd/mhP6oibMOMZN5L02U8FQeD2OIt6rjEi6geS0prNQh8l0CbiAQ
Z1M6PQzE07mg0Homcu57fSPqRwgCND5EdfVBZlAqbSdkVLP+1S71hVgpW5ud4penJ+J2jFgIqBgp
cE3nSkXlAmyaeGEzJf/td8XO2YKJA9rbQmupn0b84+tdWfvGyHNer+Mifsqcb621LoVYBc/iVTVK
aOgU5RV1FsXiLM8l2GByysdhWoNvhnUypWZgEmh26x6YAPsLmfiNARbom0wk04zmPvNUEODsGVpO
2e3LVEGbmWuwosJpxQxQBylrv5MeXI3EeCJsqouyns8E7IobjKQ3cRGTPhwOmmoxbFeeMymaJ2Hy
i/rdlQfvFt2JZJbODAzmJ8qH4W77IAyGmZ0ba6wQxsZBtQrnbzs/XWOfuFEHxWB0rQoK5vwsj6mM
3xrsvY4iqNM3G8oLZ7hAG0sVF52bneXymQc0utj2Vc6IIHEjOAsaTCeCBVMN/RnS9jaUr+PEplgq
vmAnNtMTgBFAmCjJCg4vrDAKDQ4hoFOikKs1n/cY8FocGGvls0FvEL/LmMDadUlKfA+qAO98fTe9
TEmj2YEBIrAWyOfDjZUtmW3OxwYRF7TTcI77GioFxF6QVywDkB5ebv4UjYMQcMCykaiFMUh+XNCK
YGa6wPzPDzLedNYEYeA0f39FBCTIgGOtjxVAVMo90AMKfAbSDJVLIApnAxYTxgkBDbBy3wZx9m/g
J79GIhDfDs4lIjO7dwPMUcSzjuaaAkq93Ws7zThe+JfEM/v8geUjhEI3AX140fc2cV0+1Qp8w3ze
AwYFL8pGWsEjPZR3/e9rtTaYal7ZS/c4Bvz3qtPkJsWbr+wbSjltYGt4PWiIFn1bDVM/7xksnyfY
vlXhPsvusGOWMlnXT+HV1MG7bxC97GbrN7HafnarlIAZJtjf+vIzMMpnjDcNtEji75YVqQeyOQVB
rCQxAnXLltUOpv8OpcRVj7TH/oJJ1Fg6LiX5GlrdvL02Q2xpd8+GiZAnmAxGHKm1EK/NhQQQDUut
ZLuYbOOoZlJJ1DKv7yBjEkNLaxM2p0PXrZPPpQFpbSEQk1V2kSMr4MlKUYV4oEPBjJvXE185kvkE
9OL8pxQSzl8rqOcfjSOpYHzMLhmlGgxlD9wiS/6dEZghyh//zktfoxY2iGTsv/GEayd7gkhSzUGS
E90kwHdHCVFeWGgurAPZaXIrNQ+24x/zxqAd/eaxQJ5O0aPyK5gUm8ZrvgCFb11JjTeJ6bb+9NAK
THPXuZ/X0CoiG4rFjBGyk6dIfNah2nQTt2Zq/KA1KnpbvIjtK3a8KoZkDUNpRenWwF/aqYsNcnmJ
pCcEr0MBok+0CbrJNiQpn6sJfcLl/Ubp5cRCDofRRMwA7BODi6WWPMkPvTn4A712cAI7PTx4MDyd
v327GNPQ6wDMsAfWr/w7FMVuFrxHfvvY5bV9xkuhlkP4ouV50iDRZmllsNsRLJF9Snnh5aWy8Iby
gvKBm5vO5n7BRTJNO00MZgulTF7mOtG7b9K4xj3h/+F9swRQf5bLYBP7k3+8U+1vnRx+wQ3+OeJh
7Y0NYcVZJ4lfzbezFtmf0WdCMeerKWXiiffXznqLsWJc3wVfqs55s8WLN3oq1Mb1RtpodvQseBNA
gEDBgGGs4aKdRJPIcuy/q+R2qcBOq1we3ozTYPl6FFA7CKBwRV1+GnOCilPb71uAXYras708j21C
AEQboIv2ouI0Gd/qqFhJ5oyRXm5M/qH1nYBpsdepu5iGZuUr1ivcrFFoGN/29VoXLHVWDEnQCgra
+RubJn3CmpvFi5FS2kCZbh4kJvgt5h+vt1XhSOVO9AfrCDgrCqzTh1rA5NWxzGTVHJXVyhpbuhiC
sxOwGRdZfrgPQXkh5uPkRrBbwMidR6ZHwhcdd8eKQZbKJXjHdTOhKATHnYpiGHUpOJsWl7XwUyOI
4v9BXGtbtst30V5d97h6ieHroV0+656oM2XNIH9RjSEvSrwZKVg1WwP5ekZWbamJsvyIdrzXRYi3
P1Nwz0vi4dLr+SSB0saWbmYedhkPQ+NvP43C7fAM0d/hY4cnWqLYesc1ZiiSNd+kJo+ci1TPRlZO
hOCR+HrbBP767/gMyur1irqHs7OJoAp7VNu/vB/cSI467lKgntrWSnset7FJ/gOT45RySuLPe53g
dH9t92UYwAs1cWZgvSxhRe90dittBSeZAnA81PjX9U0sV/ABKjevfj/93nq4BIx1Pc/C3QWy8Oyp
XnL/2riVRfVomkPAus1FKjFxfyeXvhxUC/lfTnTckCP1N+lBB8/6PqnxiLALF0mzecUAuHd0qmHJ
oTNmNLVPM6WJnn+RKQBiQbBuFJlSMebpHijBbONlIY+Yb7SqE9+vw5t+bOPA8S4w9MI2Xlk7AfR8
qlVDRWpY7CXeqrzXsLt4kv7IPvIvsPt4Kg7Q6jcgvg7hrkVJGlEdSX6p8d74ONoCA6m/ShT1SlAy
1aGAOAfv2M/UQC+H8jrvTTeYayYLEfNSYOgGzdU5bewrOOdBvYP6TOJcLHWYO3Ud/2OBEQeBCSYs
F/Bp0Lehed7ThAq8jhV0r5ys1xShpkaUaDuMZBaEVK7zeYe4V/lO6INik/gyIRMy5D9CeW3RJLiV
fUOY22RFaOwq8FP7L79UFi/cEneBVEYdZGPKRhL+5ggTkcZD3p2WMPgWVhLLbPiWq3OTGm8hqxou
mjb5IoNvxfPP4nIWuEgu/0g9RxpoDu3tWHwslu+fTt4IzjwfeDiDdaVEfHpOOctsZX2HJAQoyV7v
2Hwb1wgqc3LBp6wX/QWsWkR83bOTd78irTHFchABLaQYztsTKIOTri3sQhXd6WJ918y/3f9etfFI
N7Svrx5dSZ4buUS19yOd6UMyi5tC2Qp1kv3l8gja5kdq5904YBB6TRnPAR8SwNHF4nH7SdLetOUs
jzYk/a81iuBprkpN7QuFcnYmEVXW1AdHbJJZzKDupzD5gsyN1qAXyOlBf19teThkMG8kvM4HF8ya
NRglDGc8K/Z6vv0Hnr6h1mP+ANTaQn76I6r3TFV26iJuqFyCg6uoC2jVWryCWOtVEM572P0laMgj
ZihxZb9XD4vbPZwL03DYG+HrCxiNTCcxpBbRWaEAmRHIU+m/Ym2/msdmCTxIc0mZWURlFlAKJPRZ
y323+FsbccV+cCJAvPa/g7Bgu4H1iSPgXVR5PwgExSW+zCHw2rPZvhffN7D+arJ1XlBfgfW3yx67
xle0Gq/sFpfsQjKarx9MMU2nuK3sW0I7K3jhp/n0MXuFRNR6xZHS4Mq3AfUPe+CTuZrgBUqJ7Pkg
71w2B3THtaHYeXWITmI5uTCY4eBcD/pbSwY9CLqF9LcLasgmIYdOJdXCZglrHAZz839BIXX1JCxZ
36C1q0EXdcslLaRXHmP82x+sf++3YAXGD1jroNfD72wPaOJKkj371f+Nr8LvBr0Ricd4GBxLV9zl
Rai9OWXuIdFoNfcsM7MBgwlrGdi9wcKaHhpIkwqIk0JF9oKHQ0nuX8HfKEnM2dQ24/cRBpzxGllE
1sr3WS3wx7dA3fBeAvuLKOwBxi7G3aFMMagHPITNmY3RITjBR1Ckn4P72unpyrTreqH6MZ+QZK00
/stmaEefSN5x2qqDyv3guEixusuPy78PCWzbko+6jzgD8+tv3RszZKk/hsF5snlJaG4eBwjwSmKs
BbPLOJTISTEqkArAu+3/6J2Xp6UDSUBH5Uuj0bVHCiRcMSnarCpiWCsxNY8inGmKMKr70Z0GEaue
JPeURF0/waEpx5WKAvT1grjTb7Xes0pF5UcoEdTr+vdSag503gOQLvJePSeh60EbkJK5534OfgkO
x3wq8BI1zBCJrLJMquNrbDQ0RinqhPR0xvbFkeLnajvNBFc3Rhy1AFyCGZlQ/ZQoTCi1wwJYlfG6
l79h7EHVwC1HQ39ri94gk2GGFDdGcH0NxUQGSYK++BURAJzk+23cU1FxXKAC/i/wzlwb/z2TkHrP
NizVisa71U0SiUfFkztyuBEe3uFnXK4dvM5e0WNvqV+g8kLh57keF3xGGa2p+oEuWLNjeC30ZyU9
T0cKV3XCWfUcwSQpwXusKQWtXp0h4k3lpHWQyw+3s/qMUNW+mpWM2bAMYswaosp5pCQQrTamD3EH
h+mkKovCVYaTiQDMAS8cl+VjNA/6l+jLuN1tpRK2vT5MG+MurIP+Zt1NNCMTEMXBtaVzLykzMed/
3BGVlDnigjS+KNIuOroi1eTYfo1p9tpxvsliu6aDdjTvwFOIiozAAu2qgX8nSc631pQd+WjqRd/M
z3/iZsfw8zwsMW00wjBcgH09u/z1kolLsNwf2RNMoydMcRsvS4wJ8rjEaQWzlh04oPwiO4wRKU1B
aSnEKrebWcYSZHzAmnjGYGlA8gcuhE7V34DY3hgafeBbE//1uSmkPVh8QAEZxOPeXXaZPw48oHag
ZPEvpiSS8teohTvKszE8Xnv7mhowexlc7GxWuU04qifVm9BzVhIqEdq6dSiie6vKmA14Otc0sE7U
mISbcdeYaV6zjMH/fttoBW9xvAr/Bo1KbJnqAkj51EzPDIOShWP+ruaekiexH6kzRF9kLJ9whfGE
r8X71TuKTVOdAQlEdFB9ROP1KqIMTHJiFXaYJZKc6u0ojwmgp7hRcNypg1mBk+0c7SfUyrZtHTn2
eZSINHY7f2VA1OlK/anoREZX3Sqxrf5oKQCucXgTP3agv68nMQsbeSDUEf7tF9Xi7D5EzjmOW37d
/wuIQ2W7PjY063WKzw/IKEWWNNwVRT6GN53KZKCdRyORB8isK3GwSbhDIc4gpz+RXbaC6vSBEpQy
8IkEX8da/na2BjObPe1sXFhSsheBM3awQcA+1fdbdSNm2N53xfy1rBxDM4xcqdttIIBJaifBbihJ
zx29FCvbmgXHvuWt1Wp2YrLHligq9kZzebTh8jDt6rSL3+LkMhYh2HjZocWHi8cYlJYxCM/sXplV
5OtWI1yVI0bEi7wV4+/ZYyUs8zGbpweR0hmEvi6Ep/sP8+bprXwhLc8Rmx4mYwSN+ZTXuvdFF4xk
mhtmF/IkoMUCkt2ibPL3qyhuZfpnkvYRPRqJgj9YPWIBIt7fDDN4LbCtPTLy7q/l9L4eyMEj7T6S
h8gg6WfNS39hw23Y4eVfdyrREKkVEq22z6WXtwFlio/pNAJb8IOq5XmWwQOQox+JP3PKRILwh2V/
YCO7IK2/fBiVpMGuZDfl1XKKVAdZq8w/pHod32/16m6MgHXtKcmMt827tSshYvRsNlPmJaQgy+hK
MZ3iyqHYwOhAdNBVspd9OrIQ+CuD73b9v4KJTsC31MfI5c8u8ea6vR6rVUQwXyZz8fJe16B2afzS
hGsfO0G/w9fkgZzeZq3eAHOVyTGdlz8S5XA60FtzEm/b6cYRZ9mUhop2ke8/WYVJheyArPiZI9G7
xqNVZu0EREpgZIqNUktRwqIZJOGOnuA2nzoYehg2QqycevmVwwF+khE6IwNk0gfH90+GSa3WiMjO
lEqucmzR3J4xG7r/EPZhSmzCWcLENovIuzvuaGkITd1q4xaPH9j9MA2yHpNYvJYdPrTFSLvpbcnp
UmvBvnqrqJG7tfRw0t9mQGt9patp99sqafrpgN1W+vOSo6ClS/wvHknCMwvLf1HnXzDaMDOBIovn
oDKd3wzvJ3btcQGcUtj5+RcKpaoRuSZC0rpcezULtnYIJz+Vyngw8Nwg1qmlX0GDkFkKEqLesC1J
7TpvrIfbT8zOZSylA38N9BI/eNDMB9SXipe7uKMwRqDJr5MZTirteCGh4XpyNR5VNqizzghZ7pxY
XnHVIFP8ofzL2WrI0MmzZQZKFfZM7u0HLTPBin5sOFarJlyQcemlV3YcEymO9oUbrPKowcRp/wVZ
uWIvHLKphQR9jBmwHV47GXCGqXD6k+zTmNyfNOdQM3CpLG65BIFUuZBUIj1Y2Tmz7PP9RnXIADwP
HfcV9bU3UC6rFLVyK7ta6R37MJxeeXf2FjyMNskxEn0JUTM+hfpCpootGGI6fLq0X2W31evOixLJ
o955K5R/Wc0KW61ABeD1TKUOdEDi2mmRq0JjF4ixmGZdGnT9Ez0i+uL5Z6YmwJWGi/72lI9nP8tQ
Iiyd2UjNP7ytf5RILFwcBF3vLpkp0q4EAPrIPtgV7hB2FRcz/dmHMGmdQUxw9zAO14LSosLP/2Vc
L4obO7Xl8+Y6cZUrAy6U+VqFX13V1UkLU7Z985OpiBqjHJogwgiCVcb6T+EI2RNlQXnFwIokrG9x
u9ARxwHTJhO3Lfv1nViRGOzqCdxuic7lot0f2fooFf08MJhh7aNfX8GNAs2z3kvtJWTk+3AkBF7D
AeZVieFDxQaX9DsIm+caN2bLMa2e05IyzCLPHrJYB8LScY8usYmVFdVoYWO55KabgRGce/b1aK3H
24N8IxCGc6ggi56rWQlaQMu21d9TFCXfb5jLlHFHleB25Zu3wt/pKgzNQlKo5wdGZMdB+J/7XnPN
8694WsDeu8vUQDaXXttn4WkbYtn51z2qy/VVHFa5xH/otFAXFjpBwzXPE5njbmEY5pK6mKU7SFl9
z3OI+NxIaJ4e6G/eMwd9VNbO8c0B+CYNzps/UPL9h3kEvNoQZWLfZInABxzoCuLdY/vSv26C+oW1
+GJ2EkRjHq0n9V1ssc1j8ZJgfHXpkuuH+ILTbiuK36jbsM4dvHkHArB4IZqhyiHM982s6OGeDJUV
v+iWI5GUkfOzQ0g+91bNQhR26GBC84AUxYKV5Wnd733LsKiAzclrEMWvQJdevPV1tPObd/qk4tQ7
c8rg8Gf6dbrFrWMYjMDxGgiYKZXle4ne82jtJ98FUS30WlL0F3Plf60n1AgpKTVTdDcqc2ov5WKp
fBLv+bD3R63Xi4R12HNZGcFvZAXZpe2E0vBdjvhJhRLpaIO8fyYxjGAdwtjA3qicY9NNyi3t/ULg
foGxNUYIpFCPjzJTlh01gqgiBSBLZy4D29A7qiGW0nng24NvEMrqVfmhLdfEtDVx1QaKWkx28aIE
U2Xrt985/GnBPVHggiXkE43Oas9GWDujvquSghINa3kP87hVuFBs1vyjZszvcF0ivmMw0JhsE1BR
i1aGhpMxdgxHg0/gmPgeAdAvivovyf1F6yy2NMvysVp9l9jsQosPqmXmm9lsqicp0qFOThlQR/R1
lKjnxicttFEIwVboxzN1hmG2fJXoxGj2PtbEmgAXOoXuhpQsow80NuiDNXJqjIr9nmcCI3I8Pw+i
4z2gRWlnPHfcJG6PL1QVh0sJ0kHIHFwOmjiIcc8i3vKQ3TipnaeEDUX9tU0jXbCqKhRROC7D2gZs
93ZWxlmGgKk4Amd/F89IZDL7eRJxj0n3xER+pC2Ydl+BCrHXHB9xRQbKnRzK1E7IvlW5LAW76VvB
cs9iK2ANVoRyHuI6Ga9tDIjjQGP09+5aV4r4sBmnkitl5HED515DYBuYW4NSfZ5jkYNzQkVaht/9
gIGfxhs+D228hALnE4Gn72X3u4Un9dVRo9LOe/LsLE16s7vSPN8LFGbfIAs5g+7sJGHBhN41NOMk
9Kv9kQCsRNcQspdzcMZYU4Cc1CvhHpkQNvvYS8ty+AuNuUwVoZXAU9GYZ19/MQBCZAx3QFFBEF87
y2C1Ax6zkZ7XYaYi1oXwh/LSh32TKLQx5kJj+5TCoZ9EORFy6IhippjxV4hPWEVqJ4arYvIYjnPC
4Y2JRG+iswqEbCaVxR5WCWdX3NfZm5gKA4V+nLnE4yKMWKuEfksNTh9TH0n2AW6tAzoFD4RBOKYg
9hKgOgQfV6GY8gabUnJMI7XdeqdxZw4SJTmbKvTklDyoZGZnmpyNzF0U8nnWdGtFYAuitWE3hVFu
dbgVO6llHBAXOw6wQVKub91pklqRWQs89KhQpkWJra8m9wLQre/8dgovIHA1Y7QK8vVNw8EJFbkc
uzEKgrM3i8GqZgpwgC06uu+NBebXtYYZNjUL3ZfP0wfhn3QmzQxP51HrMcl2F05QJRQy1sxXQtNS
SrLK5PmY7RbpycVVr59QnUv5oLEH/BN9oUghwSlUlE3Y7LZ1RFhqABgUsbk/TfVQ7QqpY4yr+0XW
3A1nUMMQ1zPMHeJ+iX1vGoKdTbgHllcaN55t0P6fIKCstkEUxita2P2pddyY3X7RNivq+TRN3+AB
OhYLHtuQpn2tc3zbvaM9FfzOXWHg04E/ZeAB/Opjx4p33lcrcXHkpopixNDsOFc3wxgU1e9Zhvvu
iXL63a7bh0MS+WGGU34M7kP5KWO009rtI4qdsuuQ+O7fXbKSKSWlFUOVZnr3W7UdR5YfeImEL++h
x3Sfu4lfbfrSs9LRs9FVtjlEjJtSIo+IkUnMm7VUdZWOEXDW+xOZODBku0WAHAG+xlOn/wQLbMHe
R1mLx7JIAxf2IJvYYq2MhulTLmfjC5xOpvOelQkTj8l0BkSrH0grOKFiaaQp/1e99ABXLU1PmG+u
JAv6icMbh/sy/zU0fck3y9vI8x6/6cGoV9SOrtvXUzsoToJOnKUFYx2eXW8YK22PQlyNrFE0ok26
i5pihK+mK1JtAk1pydVMkiugm4RokEwgTAT3WOOmBvhck9olnetaqMmnMqU9qPaOypyn7qGcgNYq
QesAfMp1hI47Vu18Gr6bpCIRYsXRhw5hyHFbmq/R0yW7+z05QDjE/O7pc1GdnlFyF3271nOCGhIy
xcCh9bhpaL4kPcmXFjVFVkJPF4ueGXJlusAY8NR0ux9Lo6vKbmsNd67qIpSGJvcnXkwXOzD8MYMn
Yps6aAix9erdH6ZZvyYLDLMaM8qTRxzxsuo5W333D+JSqncCJC45mHGVrc0126LPx7YO/NgVvHgN
3gw59s5b2fgxG9eIEUuLhalaLDWp4nTfEClJEGdNUgGVol453Wa3MyVJnRWBuOwHRWHFmQtXGeax
uqm+SmmoLeWBIwPquvle8+L+JHuh6UkTk6BcOm2djCs/VAEMfX1LbNfSq5cQLirjgNNYmRF102x7
h6CfIZ1J8wwtabnwDqZBCqjNbchi0Tv7G640BypfoV2mn6W00fsf5yvOqbvzZojNsNbcxB8wmtDK
sBvWoGHBig0nOLD3LfbatJaYizlVF0AO8J4b31PCVerQmzfS7bhDIp/xSLuBxcIHiIDjbTZhTAr1
KSAFg4R5qFNGdu1ojBY2pOBjjmICTkvhIx+5fXLW0zRXCRm/mFwd7CGWwR4VJq29TR11Vm4VOuLR
/OMAKzyoBfnU2IhYNP7yUUo/ub+X2bhsc0lFfiVPFimWpvsWJXaQfnui+tdxMns77K0Pc02PzQYH
bqoO4Z5AdiEABkUX0HPirNqqCEgUICABJFjhOsosBdQnMkEwHkDtByrC3IGrxlrOrSidhUeWqhxK
ExTNWXfKaEpFPry2pPXPruTM/v+o1lrx0Q4N+a6IoPnVmnz/zU740ARS6FqltephuqLYRZC7KMLL
nn0ilG0oUWI+Mkz76HDuE9vQImZGG2TLcrIe2Dnit/XTYEjzSuvqhS48Yhdf0dUop87LHF43V5hA
2nmmJpSLWaoToNJYgo4gvJTbMREYcu+nJU8wf2a7iQRYmLywvh3X9KT8SxJeMwJxbXLGjNuXOsSl
i8V+iDXNwXgwNFxU0jBjXl99aJf0f//UGkZH+3XGdywYyTYL0q4n0DgQM8+9qnLg68yDVXsCzPxN
hBzbQ6mbU27mXsgtl4p4WffCeJkRP6fkSi/tPwJSov693YrrqGzorlqTIyiFsW5cq01udign9eSl
mMXVTNS4AzThXv8/VDcDD3+Pe+1siu1NlPr82AtIY17T45iod4+wGuf7/mWfdmFe3O3mchJZeW2c
NgI0lttptnztIv3wLsOoR1HBfPWDsbjpSBgkWWaO3o9Qiu96QZBAwCSOo2JPLJo2ZIIxlcwu93U9
8/9jj82UEAyBnHeeyY0J+Py0XpTaOMhrAbyHyqsR1ZlcE2ALldQ6i3vQ4Ts2cyedhzYPSSqbji7E
jIdMyxkOZd1jpbvyihqplF4tyICq+sd8jbaujPE8dGHOsNTY2kIlOwzq63sgT1ADH29m4/fUxvp1
1+DE+zue8XWr3tnW7KKU/XqvVKb77IL+OSWUhgIpfYIFcWPs3CEUyWrod4cz79m7loozrq295FNk
Z/ulpKULx1mQKiZOuKGZzaESbifqBFWpqhhtFP5emsBGdvLPFdHrolae6IXMGHNBJJmUEOolw+MC
HxoN6P6L7tij12mXhxgIm6Jrg1UMsO32Jmw6uT5gPTjWkcdpk+99MYhVoaUeBOJ5ewfxzybqIqYh
XChgK1nHH+FEe3vhOEO4Ufw0ZhC+pF73PxWGNRqMO5NVQ7TRgyPBsPR8zIneTcT/IvhJgpLAuHio
3UEkg8v8/iU0OAyqEFczetauLwhRKDnKTS5pKdjpZT2RAlg7WrmtlIV/aY1gYjFerjeEa0TCKYxN
I4tKpWn89J+PIpO9Wc8yHvWSXTQtOmKPD6jVXPHpWl3wQlgW0RAuG+DPXBnoZapu82bN+n9XlcON
drGqpcc39Y7ewhjveZ4RA1lGwkOfQC8kF0b6SqNPl5Ky8YAr2vIbNCyjjoUX4/Lzs20xEvbZ4tj5
DbbWXl74U+WJUVCbovY0ru05YXzAVEr1degsYqdlycSNq9YEJqG+Fkj4zPp3gqXo4xnj007KB8ai
6yYMsKheoa3y6nlYvGEbolG7kQRPeRgWGZ81xD0a3K3gDI3vB2qbHxVeqSlO39dK5wCgLWc/2/B6
sCmfnBnPUO1XyQMxezlqsGLXURWl/KHZejiLQF8DLi848Jfw15r4DiY901bgcsmo+ZybfNqhdfhB
o9fxpyB8YC9Nk3EqQVSnJZUMfhuxhOWQHy+NP2+v7HypGCIgge3qhsBNa8nFOTIpFcw1tnfGUIXD
ydeb8HmwbIt2vjKCEzlOfsCFJlSeU99j5YninpF0Ctnb+6RZSxXqDtHX495VLl6HYENoI/c1XV4Z
4POBjCBmfjdfzMUusA0hrx/RZ0kuZBL2hbs7CvjcFpntxBrNwuYMo6N/Q5pxwbgY8rDbLkJjfN7J
KwI3EegTeoXiKjJRu6iVykfra5Vn8pFq4EfxhmMVgC23OaTBvOGJ49mAoXMEYbuFY9hU8aiieior
gmITaSdPXtKcZMIPXNCDw/rYAEYajsjWzVIs7I+fL3yPid74zqXpkcaoAxW1qCcUbye1cY4ttx4A
qOHRL1VhnPizP0eFYWUGdlL1m+dVXy2o/wtyN8s04DN/a3+Y3EAiO6uS6ba5NI2Zgw92tDlCg4N/
DNmdvCOletgIh2CEB7BjrxPm+P5G2rvyKa1byKVcuEjeBBTJvZTYHvZ1PKKouUYGKe68IFLXiqIB
snlxo8pwfid38glrtx0tFN3ExY6S3qGDHEI2TW3JKdUOocFYH9ojIURXEAZOVOcbJQdSumWBDet2
BJZI1cnD8Pk3DGUCxflEp71AsgjsruvpwLvZMC+E+mdLJSkkZutUiCx6DXaJw16ma2zkubFz0t3C
D/uEXEWIlWQleUJu3mFe/+r2h4V5a7erK9ImWdmRKVqXRdXe4nnfp0znA7rX+KWFEA6ICGllUY2u
ncw1Jedh+JUdDUvsxzcW8MWZaKg9feSz/RGZQdLdqS0Updgcu3NiZ7r6IDJ0THQ2xqyXKmUvhx3b
Rj7lgaEVpjoZ1mF/54/P13x2nXCBo+hA/IFshYg4OxsPtHkgWmSAdMX+4DKUOOMo9KG2maWHQSnP
5W/8DyuvCx/SLAThxw2p1Ff/zUUeeyHxLN1u81GGjqqZ3b7QxaIxvHUA7ucIbxQYpC+Ru7ps+Xs3
pKdAiiTUoxgZOnNzhW1Z/41XIhxaErV6MyRm51sp3z6vurrlZjFvfWRhb1xrZ1nUsNSiqkFHkcyA
2M4wNWp7PtyOnIdpYwMy866/YC91pxmVfuHz6+Q1vVhj3XBkl7jPdKcNIAFdMhZsJEPShWWWH0Cu
usLiG1eNdOKGOhEEHOtNnY4hpWC3gGcounysLvhqfoeAAG8zZ/LUJs2hET1ntu7/Bfw6cyv68gtD
TTgaYTrV0xKHDoNJvhRhc/8JiYZsSggjO7gnhJa0RZl8q6yR44z7EoY8izseMhVLG+0OFPde7L0Y
9cSfUOxLP3a/p5DlBxiuLf7VpPgR7iiHjOpHpqiExfwrQ7I2RGAVcs/Lnd1TalfztBM6O4ZpnKdm
4uFkXsg4ZkyZ53grv3/eFwqk/bzKqwQ6u6lC65ctRwlCWrbeKSfkDAeWKxDzSyFpsliU8Px0SUDN
TSPukDQkh1Vw4eUXMCDlSdGsl6UTW/1BakwieKN0q9+oHHwrzvglVm3J0/wBOm1Bfx+ih+Mo9RKB
GKYov3KQXEF5VmoPzZfaaFzbeyJzQov1XjXCl40TuczvSavn6pz+sOc+JNwzmwMxoD2wSGPFh4SB
PpX2PgDfdp2FWKtjy+WhyzGfmbFw3AwY+Eu+kRSaiExXkYis0H+LJWEHO5BCbSrjMquE2rCSeirQ
09OGjxaNH6Dvb7d+6LdFu0wrNRuVLNgbGpw/+XdOWP4K01/HGhXd6HPOxqhQtdUeQXl7N2R5kk1Y
MbREvoI6gyt6EzA/iMoOMlTF7qjdm0IMtvawnF78uLQcn+lBwi1xFQh0fgQcpWY0j98/xEfGXH+o
+y9OcEYxguTAdoLIgkRL8DQ6SIObHKzhBl/B5H9MNnUAPZt2q2qT83tqhlwocDlpUI8gqrNADo9i
CtFch2RDrOWY+FqwbNKNgBExjGAFQGyEsNCyiDoJAg2DCKhTGoBYrdOPkdlUIZtOimvBzal1cLLl
Im/hZM70TITDxppvLE9X1j/3wSlyeRfsNhXufcGBD9hcG9CnMf2+KCUoAyqYigVCxdRC6VBsDwpp
1pQ9qw7r9BaMMYzclpQz6y0cGUa0TQIZWiQYd5QECVfO/r9CNlDfHTMRu3LEZ1v8WwM7g6Tubki6
l7kCHeszEySb8llyV6ETMWJolq9nUR5krenLcNDkKNp8MTI+/dNF4yAx1liEyF9NmrTJXCyNlAU1
v/U/xiBnOF2VDoWrUTDYupGS/bhRerhRDm7cpwtdBjTicJGhtSP5ebD0nCEjvvpp29tcaK0cEoWm
vtkVEcp+tsSxQn3PkCncmCCtLgwgY8YkWsn+RTvRc+6CbTa/GRWfHiniqt/d0vscgLOZ3n8+yivc
TRff/OcaoBtltdg1hjI31h++Emr1lTSzSHKhByj3LvuB3URH3tCtkgZ8zRy9GAHtFU15iO8JbO1C
ipqqnph92gL8O9TWX40NHgYDDBivRLWAUEiMZgLvTurxL3ijxgPu5z4mxq83dOnEvNDXy9p3BnKT
Sv73hiXqyrCVPZA6EWVlNoZYhQufKWLRcDyA6jdII85ZG+gQcN9keTon/imhhzruA+GwO7DJ6egc
9O6pA4aUZ7DMsk8gB46ndb4jzPVLAxnywUfTI+T6MAYVYF88a5I3+h74yMj4NHusHrtVweWGvLj9
hewi+aaIFvpawEW5epOKR4kMDbemSMJ+M6NByfGDfOO+ll0MhiYy6rZHcIi+lrF7cviWBIdP+WaB
+pB1Ry7XiL+5rDvmb1rkQJLwhE3p03NkH3Sp+OgWqVq1R7ym0mZjYleo7WWjp8pj1wWjdYZSIs9o
GD1IuHz6/La2Z6djqvtQZgDdadhAk895+fIHMCdMlWzav7AUDrYfFrDX/EEzCcHvHqTNPvgFbeit
SceUcylQoQkHNLhsg7vn9PhnnhnjYCrn7eWp6CpyQ3UDEAB5SW/3AKr7K7QWqTDQ4RQrU5KJ8rYi
aJVj0finnpZeWjLqSHOGq84it90fS8nhh/9pGhG9tMGPjp2iIxKvdo9MysWJTudzbpwzStYXu7ZO
KDhWYO3gn3CsnZ/2tti1xUfDu/KKws70yMXDNasnV13+i2u8ym406tGphT+4DWrUizj/nYIDNszU
5kFSrVYUMEjjwwLx9UebxxD/QzkO5FYRI2E9AB4iMGnIRFe7HIEIljy4N1MYFl+nUwZZf7F8Wh30
sh1vPaSspbRdr7CX1jaTEy0TwU4Bk0C528hRXmTi/pi2kfIX+T7McvZrZLfcK+ZRHP+RVi8fBY2u
8uDJW/Jd/uZi7wKHZIzaCQxPz4FgS0PBPmRkkxkS4tWGzfqHCny2pCXhFP4CbJpx2ZicdjJGef32
y3UBWUloOVzQg9HseIETJNmjWmbB0OYcRAhiwi37EuI0JYorQXQZk9flI0GMh11OzycbKYUBUAWa
bCidRoXpLAtZ6dxssfQWF4PkOiWcq93BA27uDaPw9b/mIPL7HbP6ZOhjF9ribNlZjA882wvzVAUN
A6bfRX5qbFndFYBsXGHkJPCnx/xZSFx7WWCmfzOuFWJ3IgGNoZrHWyVcjUnPY7m/Vubp8uUAp+yB
+UYHNScHPNvRKuSDHcmhWqYGKBmGevOxSYyCj6aehInGC8Hrm+thYC8r4jd5Muqi9r15G75jVmAP
9GduDJdazjQ2/CUIMrMg70F52JqU3yFBTwnX7L9n4G4SU+ipfrHIQU9hM7OWSyALcXn4qCjBRoyz
BtRtb3S4UaYddpPeLafAN8st9ISsSkSMsq8QR3+FI/2iYKIGP0+jQZ1A+pBtUC+ggdjKrOtic/RA
5dAEFfCw6GlD6rLXtv/gxa2ygklTnZffhQXjOlmNBzNaJ7qcBIsVUND5DbXiqRQJE51FjwrQAmAa
2D9F0wndEirNzLdsmecefHYzvpjcmoWU/emRF9R5cDc8LFXzO/N9d2mbhoozc0JnUdIRd69KETms
P20yX2ZZDj2wqsEFEWTRH2UTI07n8oyFlTAhk90prxpQC8PWBUViLDpA7p8Ym7w44EM04d1ERoTN
sFBb78Ec5U8rmEh2RUw1C+VZ/md2u1kzZsu8oTM1Z6FccOqvzaY1D8/EZytjLtfWpFDZLm3L0IIN
e00WfdoxrdQV8UyGYFXd6DsuiwOm5MDKyZ/tQ7ja6DtZDgvoeNQaw0vSVt7b97nPPb8bnMWhnKrF
tm3PKfEq4Fg+V4vC9zNkS3OxfbGdTcBYeshcnwA/47XHqeRHP5iM6klit30T2XqGvtq+WAKviBFb
Y/fCeQQSlJwYPxzcNLzMyNg9e6zFKn25l/iNoYThr+HLNo+25xF7IHzQ9cspipDYgo/2iEqNxRJ2
v1UAdMAODeZKdohUvJ0oTCgaYOl/GSoCo4oxMon3aIHEXEafnRd/p2Z0czyJKrEr1o++05RE6b28
t96d6oCjvPw56WPuCWzI68OYES9NDrMRL6nrZXoOSFe+siKWMRmDq3FYzJHRPFCK+PJ+512fPqQI
d5rEVIiOetmSu7S7FOBvvjV20Kdi0SR6pLsJ/myexa59wWfZvBGtQFE9pyurl/Y7Q3Ii3qKHAiKj
kDQmd95RKRze4RUayHDceVgrJpT0Tgu1XM/IGVmhKJPeuY4ruHm0cO1sndzs2vqW7FKPEN1jQ168
NL2Mbn+0ExOWlDDXRXRbT87SEGsOCHEuW5ywc5URoC+v+baIje0mjENAe9wfHTRMQhHJ40G6M3IF
d+Umw3VOSp0Z4fb5nJw5ZODILevTg24BV6+ZjTYeyd0+FQfdAXbSJ8T1cvGLhw19K1P7+uV26go9
zmNpuu+lqlfaNAEwq3hCHfwKriaKJWjxpItBo/PhxW75+HjCuLkQCR7EsbA92C9rwA+Bv1+zqThe
eVGu/H9B65Oh9icjthe5Shmm947F0gvAA5QZgyTzIdlShgkJB3UE5txWkni1zIQSTxLFSkuKcoaG
fhtRQFI6w7fbcaHYitf9wc+D91+pgzXCVbksXiPhUPP+BEVzJ6UrvGLvLI7tra3hsiu943kLgkHH
KDkxgXgXWF3XOAlqkaXA8j9kveoaMkT3H2wjcxP2NC209CdhCpxLa6yRj2xuhZ0feWe7tAcir06H
zm71nOusp9NErl8fyv7FlDUIliytVNeqIuNodL2AymFET4EungRdNlTEFZzyMXXmm8LaODH7aeze
lLA4RgCCFpwDl5EcKeYRPig/7pK/sXVRXjMpcal/9YLTNa+o1rTJHkJQ2KKXYXr/hazr7NLpK9+p
NRv2q20yJAuqBr8eS+o0/LLMTjj7lTNOLuLXVmfwyMjSgj32vmgVac9p1Wi7en4jlrJv6c66wUMC
s+zbRsGStSmsQZ7R5WW1Eb/VbOkCGqLd+hIOalr/IPQCWSDFoJ/Lsg4DcrQ+CEEHyGw3T0k1Vb1G
CDqBEknHoRdkUF4eArRWhmWg2aO2b0PeZV3lW895W636xlTOq8VxqU2owMC4kF3jCzKEHIPYKBPf
HLkDQjzp7ObkucpLQ5PNiI0q3dA5iKw2lcCNDBqy5zOEYOjgmdt2hiNdU/30WK1tAiU7YS8k7pv+
rdJOP+Gtl/GliJBX8CX3+dd+7YNvXo1Cw6KySO9c7HRuiN/V3epU9ufomUox8M09NKjI7dDUQaNE
QT9S1C7T0XjHOD/i4szsSSn8UhwueoNvmrhthBpbMAkHMGoJBL0iyMdeRwL0PIPFbX4kbrnu93UX
362U0F8l7SgODQnZcW0sC0AkOV1Nj9LqvMpoM5Ssxr8gC9ZcbJ9qFH8t5eTo35pmeZbLGtxqXPzV
LP62GD8Jv+hpzKocsi7jWfkPoibHm9/KFISf4COIAr9EqmHSr6imE7tF3wQFQUcAE4wt3E2naS0p
rJfNoMmTcAbC1FeL6SGqyRtfv8NRaA1c4UNEBnRpRKpLY6pECZreEnP7gJft6s5+qeMZ/uCmqf1Z
GWQHUo45YhF8JjL6TEYtK20B1qhAnhZFd/FARM6WVIXrrv316Y59BzCxh1PQRWsN5KwikAufcbc4
SNXIUU4H6vxuhE8vkRilKIDgZhXpoqamj4rxEnmrBO9pMT61aZMzanUmElQktnH1WRPaafOxfflq
jjRixah3fFch6rgW1yXgtcNgCjoOFODQi0YN63rxhCWFJhXBZookZspctH4HditraHcbjCCVzNNM
ZO+QFt3qtx3HOE8qPz9jT3a76+LZozFJI3/eMJkZELdhe8nRlS43ntJXfFWerarBC73G1VXc6H2t
X6RaaPF7NhlOClkhaCcw1Lh5Rdr3HpKDmgb6uQSnO7XpEU8e3G9ByYd+IdP1gZ/orrcdiLloqNIz
/qJbO9vUmAs5KolMdA68oTk+UPVWEHwfKEvWJ0yKY799Dl1VdplDvRmoN+a8oxThsmFneIv6/YdT
oFzc63c7OGnrGYS029SZOZpWz1TMlkCz9FdmZCPGtS7UEDFO1pmlucvtdvFLNWnkangyyXV0Audj
VMmFvu5fSmtjk9v03B+wWKoCBO8zvqptFaQS/CPymxXdrzYPAPFqVr3CQvj3oHTDT1UfPqPd1Q5N
tVpWjrYiqLrYQOAS6BB/bUZgJvNczURea0WyCrdV4xk8bOL2/RMgt3sf/8Cx07hO6/xnQx8sFvde
xCZZmRF8htJtAuMSltomltbBcAwG0jrpwXHh6ODS1HM4/hvcAP44FdgCIW8mgPtrf97ZeMnDIU3g
VNd7nKX1w9KioV84N9u4FpgL9VZ1WGdcdJ7IMGpykKaRRdqIVc4LZtscSTrjaRhL78EKGSQG1ogg
V8jHKMdzmbCKyALmt0lh8AZhcN0d9VAF7CKYNNLK2g6ZFNcNndYfbpBhT31uaXeJBM5gU1OyzBsH
2CNkMRfvekuEY3BYrFa+IDMZ4GmQHAEVAl7AqZY1iP2akSUy1KCQtu+OtDvfCcIrUqc/0udKlJHg
z/hgS7kQU7bb94Q1SZPm1dd1AKfT/eBdkxVOlP1RD9aty4V10by/SmH0w8Rim3GRyftZnCBcI50h
QsEQqDn1dpGcli1lXE9RFd5tN96H47YzUF0ID2d5nH4lqZiy3RqnbueIf9+pgKcsy82g0Z6VJFOJ
pEKMqfuq4rK4rGEyg+H5qyXuoxIpymiFyGVLoBLGxQL5BkgcGejb9rJLq9HWvCO1P5TZ8tTRv1kc
Vu1P64KMm+eN8iBY9tuTAGsZPgFpHHaNKZsVOZUVhLWF5OS2hjcv2RN+RVDrosD2T7stVksYeQ+v
6rnmt7uRrnAtZhV+Bi3sl3In29Z9o40xU/Nq4d5RuWU/P+vhpUyldc+OIE+twrDWt6jTZp5N8XJq
Jbx18ZA8gKF6v04+ozQDqcWe14443yt7DeI3+yQLtiWECQGwAqrpSCbK0+JwRQcPD58bTx3SKPFI
c/hbpCNSTGYgOtixjaPd5yDzSjeWRElsVtH4IakJ3VBs4+QAI3wSuxiMOKtUrE5AMRyMK+37Ob1T
NkH7pzaresJ2scV8WryJaXkWv4fRyoL+3fLcrMlg1lOUbCVJzIsSOaiDnj/WYyAvVPdV9TayLMJr
+3N1p/DYElyqj9z7fn3L8V2NuaYhj9pxhWGqCJKzt/D7F3v/JFF/zVJ2vpeP6JfEjy7pXnCd5LsU
A9an6Bto8Ibl8jqjoUnjUW4W9fNyTgKwwjVhiMsx4oXijE/nYy+Lh0MqZDlzfANyBRkzzdOpkWqQ
U25dKi4YFDOkZ4IYIklz78AQGgUHZaM9gr3hMB7NCfbnKIwv7/KwvKvJTOxstC2pKiEgTtZzm/tW
s/ekfeDZ0CU/Gj2PgrVr8Wf4gRtU1ca5c+Cjc1at8GR7AVAh7siiNxf9ZxDD3YdyQCbMUUPh9ugA
TIcIna3Hlkl16Q4HGcHY8OZqS0cNNo/h+TD4l/cbPp1hMdqKFIQavFsyCnKJhYtkny42roX+8KCX
AwCNuQ4L4CwA6WHwt9WyB6k3fLdooevtapT2Vs5G2zF3DQBpK3/aDpiUCz7m8aoot3xGLFmxSBfz
c5eojqOUio0KREfU4h02jKDfc0u2R98vJGHADZWMhjmPOty5LWreeuUpI6M/ijL5p9nAfDa6337w
/ie7vlhtzzJOEer7LtloXzTRfimFS3e6CMdOhp4LJvrJb6tsPQ9QkIRNU91mkCVj0d6gTd/rrUlf
7U7mbc5l4EKQ8eDIHhmRDngHb6R5tGFlP1L6lCKxPA1FnhcFFl60WIpWpEuKeSZHkyZMxuaMkwHU
Mqy2tNo3yNkfOeC4PNNcBUFe/cnIbSL/vfeu587zc6G2D1bnm8NUBIEiy8Mm2UylvX8Cq7cbZC4W
gg6jGQ4ajHSXWehfmCLlS3OrwrW6nHSyeau7vw/YnflaUZmVnyoPM0GRyr8LU3vft6sYu2zU3mJl
WGT57jsRbD0oYq2QtiDw9yoGzpGBL7Poy7dnRjBcqyM2xSb7+3bDG3RGYwgossNwX+QtVh5nLF9j
VWNTRs4yX0pIQQlxwRKHYDbhleTzuf4GACNCwrR29jLm2YC5l6Hf9dK26VwIxIOBNwL8v1hNGWf4
p/fXGqbHCD4F6GLmaD6cPSv3D18kcwzFn6+s7OmDxrl6hwxs46QDdiHttJe/f2GurbQ8qG6bvisN
jaggvViLg/K7yAIoXfV2ZyKoI9LH+DTpGQT7QebTs3/EdDvYdsB5Yn1b1UMPMT6L2sEBTRf0g2ua
9/L/H540XG47w2uGmj/OVbzqRCHCPQLelCgGR/1fiEZea71X2QW9FZ1xMLxVcVG8oG9PRxMojKY3
Htnv/JF4pqp6V5zQJSMJxHTRDpt7oD2Ym3XuQJoB1x1W4Hg4bkJGQzUFtOT3F/reGVk4RdRUvHFh
ZkRN1qMcGnL8G5m0Is2Ppqal+0sP9uNtK7PG3sk4WFG3BjCpgA9eVJH6l4wMC8/ooYYbmZzPEiz0
dDYI1nlvWqkRRzaQ/h3Q7Tztvv6ex7a/mo0cDjvRaOlMKqDkimDoleU27RRWJr4UkK+k9y8VBrCa
BzWvSzPPa23oj/YymDXQZ8d2s6Q3M3FhaAel0OAwUw8EguorubqqxL+xHvZd3ymfHZy6erzJfEj2
31rCdTXmqZsxid1ENwUnPg2VxRRwl6RTdg1z8WTKJAu3ZO2GNGeT6RS+lqDV1L7ZDzux/agp87GA
K1z5DHTPqf/lukFDkIIz4GWqJoJ38ajLjt3hh2Rcg8kn1HOD5Owni9v/z18rLx2kFilzsBakLeCg
RiRMRg5p30+rwkkpL+nWQBqp7Aya1EWRWNQtjUrPD3RBh8iB6AyLgBCqFuodnenlNhr6mh4wyEcM
ZW3PfK10ILTLrpL8AXjYsPtU5Di0QJXwcMSSnCV6EoV4DBpd90/iHBEA/b3xLGkSgQNYmCxtabw0
LndcZua+MvhtItaNeWqZIzSHtwnFf92c5uXr1EQIf9Xwm1+k5dGg4gY21h7kDDNHqiUL0OV/Wq5r
7ruWJ1US5Nj5oWS/ujRM4W3bvH5PleECHzOasaCHCTu82jDeea6dVBHzH+mwmFHg7xbXNNY1GY7W
nSphbrmB4XMCjT9jDsWRpdbbnx2v7esbL3CbRIPjNdC0xgMf4OmSJvAJq0qVhU6AKmjD/Yz6kyo7
SnaBJ/gO1OpGOwwke39oImZx3ZNOnM4YK8mbFv1TlmTSV4Ko0j31QX7wHHACY/JabEVrCFLKG9m7
y+yMIz77FiGpLAjlkau7nDLYKwbn/Umbprk9VCywuYaWOBlcAST3I8Wp5PX+g2X4XKsurNC2uN6u
jUWR7bqyPnq2vHHbC6k34+STQcSQALGDVMaLu9TRQc/R43ApW4ZKHr53AQdI24UXqdxH9bNoxlz2
PVTIVOqJX33clYqTjf1BTqJM3TbzzwoUsKAVuQ+Tam1k9zfyqA1il3Unmdi4Y6lmjyrkjII4s4xO
LNoF5Zrhnbtdcei7v9ZqncX43GqAA0TrJegc9G0IHREKkYOHKAOu7FAEohSF9vyGWLLzoTO1EOpx
Cu2iYxNfszH7CZ/ij3KVTyT5rIXmPosP47cmxbKPjCG4ql6Bdq9MmnFHlRo6ufYcR1eLl6EcawGE
Rpu1Ny4dHXB4skFZzPZoq6Uuq65RUugrvB8NStDT3Tce2pr9U84sNcY6EaxWA/r87iU8VDfj8I0s
CJhDV7TlDsfmifSxRZVMNyxwL8J75FagjJLl43eKXhBxuKwIa+DvOQRQv5EDYmPzp7gV5FUBz/jq
Z9PaEtFChF3wisXpLHXVuEYAzV3hVzKU0mWhJ+rkAtXYLMaQMpO0Js9FYfhIMjCOypQuh8h9HOkO
oDaceHdn27DRef9STZ405wgFBhVGWx6JoBVfnCk9oG/8wR79IeeWbKfqupDgRzOBGOLlhXVUg0jF
r8AEvEck13UjCvmAAg5BrrsraXUU3SpQJ444iZHgncx7mT/NHggRkp2ty5KUa/eVIk3Asxzn1W0+
Iw/vZI476CJoh13kTHa+PV2FdgeDp93GWBXPzBSGvEDhLNM9zrxG4kD/F/0fxoRTijL9p4cUyBnr
SXFNsidPU7qANbBfoRV1axrdAkEhry/lzkSTLSKZAq2QdgEIVqwGD15RNEydytmN05MLMO9MYpd9
PG/JoI0leq9VUjANCd1OxolajOb4YD+aQKucl6BTXElr4Nz4+TSQZcuZU1mYlYDKV+ctD5Pszr4S
gelG4u2CUwQzzfMCfVR8Dpu4HOPPV7AwYS5YEfMK2tCiOqzrJmE/+XMPjrZTUPTc8fB0+VDUfV5C
l88U6HMlDv6yNlDJeXov5B8Vmkxc2b+RAG7KRpUqxVNPjcXIZR29ycZ1IpzGEe2sdjQBegqpR0fK
ekQLJZifbJe9GJLcDawl3zU+Zlqlz5XblqyIXkeB2/9GMFIiXRgXB7P7ebVf6Z2RpvIeFffU9kgU
9BGOxEx9qrt5f7avBWtc/YCtl9qIsRSCEQgekjF4jORs0w3EiqTdj8FcK/K+TeL+nCvM4Y03QdqG
iDCfJSFDhTOPfDT+Ydbq0xHqBYMaypHoxUCzaBuQgPQeqZVPp+FKTsQACAt6GCBN3Bk4D6Nwxq+C
iJxeVv4RC7DhPvn8ASzUMc2k26iU60v7zUdefKIcJ74IrvkihUo/c3zUb6Ta5RjzP7ZRbt2wtBFt
/AdmfqzA7J0GeKO6wOe7afK7NWQAws/vAcu6vOVcAKAE68RBODPc64o8DPP+hum2nOaqF+oS0wEp
emSIlmuaBuM9G51nzYvpg5C5nXgIUR1Gf6XU3T/mz1rfd3kfPN8WJY5QCL6zHRh5nZmWPS5EP+/h
QXdIHQqL4CLtHXdacWfqVp/h13aME8FBUfCMkqPDmTpDDaqPZdJzMl9WVlgDMm0Q37luWscdkRXm
RbtNjzLgTHrYSKhE60iGvxcaO1DqqTO97Lp3gCMh+H3tf9y4EbSlsMdzq66pj19v8R9CBtzvHuCp
X9e29Cnwk94u3iUlrXhBnNvrikbBaZE+wjdcpNoY66SfaoRH0OJHXIAWRYCQOpEyKbTWKRGQYqFk
a6KUDqVEXoT+5LQZz1eT0pijLy4//11OUTRAy5xB2ZeAy2SkrF4eNaslMTIU2qhNmn7/JSL7bqC0
+6V3YM4mraXZuoI2VVVhQPX8wD8CaMLXxEvCTqilbn9i1H65XhvfwfHww2lRN2Er1V/lS+xdUetv
ETOCPIzRM5onktpsd6ZmpDQQlcLi1WIg+ZCdO6+g5y7+8tKRRZ1cGTXWYekhVni/ms8o8/rzmTRd
WtLv5qrJzTDD88h3WoimMri3XubqHvIFo0h8+h66OuERUhJeewSgbxdO6OD4AIQfyfwrximeQ1RI
KZCMVnsG5nfgHRITVLkWNmGwl+sXT1HpPWSTHpiYJIDalG8YHav2Z243yTmZLfO7Q4zI5VqLfPun
t8GXnoS0kTYftpfyZPol6uNz2q+6K0+RIjtXPLABB7w943iT0I15eiGhv5KNUA87DDzLq4GeDtCY
rOKfKZxwWwzhMrbhdjG2UlR+HNL3QFKeIuJ2sTnhHjhEqESdwUAeeYdeaW4dPzEbkj/AReiQsTO6
1iMtZ31MVSJXQE+QFzlGtayB8sK775omSlk6EhU0bwKSJWCTTfm/pSNuaCjTFnqFSrMOFGUSfaRx
IfXKakIiyzoG6i4p2Y5JomD6euEVTw6CLO+zAmzj9QMzeHdC71Q/utXpHwJE/bbkppU5Vk57WjUO
mGmRuMRw4LegP8GR/zm4wv0pa0wv/Vx5jRnxMvnSssNKiOxeSR1FLxA6XjoeMsQWgG65+eVm2n2T
Wloj5UdCs6eo5FWSHNueCGAnejsVMIHpAOayHjJHp92qKYp2Mv1oxQ/D9uPESgt9uvDHZoprB/n5
GBoWFMnULrsTDoZho+ZKxlX1wRHl97LoF+QYP/NFOd9w8MFa7ksqys9fdekZ793XnQ4IPWe1r42Z
sWROl5LkZ5jZ38xSijKcA0r80T68qGWaUYKO8BA5GLDtfAZDuKd5ImcEw70kQLmYDJHTOM9ppPRK
9ha9lwuD80/sHViG8ju45op16Ick+vK6VWEtXVi1qdgB0JvbDbxnChnGulFzAHjjcvHeJ5uKPpeR
EfjJJDWbJCEHxbS+kA7zYmhfRtOQTtXLFgBQBsnqV0mWMg1ovvxNn15pnUgsHg6wBdvZW/cLGCOB
8TVxboNQNABj6EZJT3rDwBFqNTG7FY8BFTDLCIVjN4b8MzRINOURfHrwpGPTrOXcmEpqzlrvv0D5
AyoTgncdCbIKWaw3OygPM7Zow/r+JnPcyXIiuAShSlbtUX7f/qrvgXaxBi3X33OXfh9ji5Z050Qg
zUH44ogXcCsf7Rrte07hc37ysLID5lfkVrvjv+fQ4kT144i7tcqorSoNo8/7IWtLVEiqTCkqsM6i
xNfxhZcpkUN3Wn5OkLtKkKBoji3UBcM6GTeSnwxT/lEVsC9auEiLrDRDYOaj4jMb8fNaVCFB3bsI
JaErdqulUdRQPSTH5SlgEIKg78liGsQ9BMQkdzpOgM8IdKYteWqNRhVhg8+EnerkhRkPuRcuFyit
VWAYZCcxKbyq7osZd6V69uyOkx9PE31NCFExRARCu95OrbdPrlZyQSUzvQtAshX/sHAMBm1flRhk
sExHjAjXq9mitSzETl+BsQFEyxi0OwR59zWoF8Aph9/dF74AcPjz7ehBE25Y+4bRUoC1mlHxHvjD
kOwXOyfHW+M0ghwhWwSH6XI1MRSFIrMXsiCBDtJqtgFENdwNGlmXDVfkvWAWMOGqhD3Hn7JqJHg+
aPJnLOV0hEnPBgMTj+VOO31Cs6kRcKEovbERSSruU95NRKY9K8zJ+im7bFDgWqcCxtNTI/AFNU7v
JXVDK5M4mEpedL7lvym4xlhq2toDMVZ2aL4BbC4nMZN2xdbVwLGQfCUHIUZH8XmAchMlXvK8Zuf4
8Scv+jGQEc555Z59GSZGbkSGWPF3hSdjmlwtirU7XzBIjB/BXR5xOPiAE0xAlpyvRgXkAUB4mWy6
93TWDyI3VQGAFb79eEMsxiMOiGWYuvMXoTdJ14UKssuOGdzJm0E1M9YZ6auQkt11OmHYByfZZoKd
sx8zraVU59M3l6QeMApALtSqhRpH6d1Q4d5EWygGvXwet1HwVSOz9TptsHpDCDrdNPA9db3N+wrG
ekqJC2zMat/NiDkMw3TFtDOZSvIMmNaTFi9qVLkP9N2ZSrux3wNebnyo/V5XFxiw8c/wJo3DZD2D
rspzM/mdIssjnImgCJVkhFsCX6zsNu0uqN0WRuv1c9U/OGy9ObNUWLkuuMjv6Qo4ziYKP+acO2/q
2mGKds94JKy9JmJPa6m408N7LIpwCQFs5hvOOEAL1+D6jb9kkwhBCJCLxKucqaKNwnFaw+rdb6wV
PmBl3+pyPuiwMjxh/ceRS8MsXcnnATXbFHdeVOb0iaBw287qMRcqxJ4N7dEPDN3MmjOF7MsvWbLm
XhKY7iCGNt9lR6iU7Eg3w8S33E/QucL69mEQmWiQmoPhAhiA1Mj99At5zClNf7X7EcSd0VyZqr4p
tMI/tmFZwZMsw0CuXhmxSeYsUoOz0y7UWlkKlDIkCDArMnpxCuUcltFyGKkC2J+JB9hLRy/oGo8Z
s94+0iqvnp/xhsPyiWZ2gjl0iveucFndsOMtHJhBwXCGHluZJDgfxXY//zG9uJXmmph4I6+uvrP6
7GHX93so6KhRKuJjYmWghb2ih3+IW3TFXzSalwAvzhMmwVf9e4g0LjCZfoAWJLeKqPauMc1ik1rs
7KpyGlbqqUVRKy/VRuyn9ZJf3QW54Gwj05ETMVAVTeEe0TzxazUOGHP6/3lik+W+vnnpU3jlT0n2
l/DF5Ghm1J/oXgPoZ72PUy93zmT7y0VoPQaXJje6u3lDapkZH+4L46PWs8jerXk0ebreGUs33G18
ICD4P2IEuReIJCoIHENtLNXX5eGzl70SB3Oj1kKMnOH+Dc9D8/3xaTHrQYvhKV1oe5QVxf46zEUE
JTD555q+ZqLNtg6aAMw4KIU8dItjht0qAmUcCPWiiiDh/SLmNzwf62o1nWq+cPLrZMrM2mM/gDS9
GRivbcgFwiRpWPFEZ3aku5Z92zEhG9RT8DlV9/C8CaBFwW61t+li4A9Rb4DWumFI/7NCRWUuPXio
ufdIeDnGQQV1aI7R9aq5kifKOotWHpHzhtDsxZWhnZl68H2hjqpZ4W4njDaAlkGMY7E+6PRAJGUp
I2T4+hT1Hm4c4kjh9mf2nXstJFJMMt3foozbhDLadJV7CBqZ63h4FEcki5cJPd+RxeoTX95cxvJP
T+Kde6GXGkY8Lq+NuLUg+QyoVplM3ZfgUXL/2X5uDABhV4mvovAR/wMmPpbSm0qiiyfG8YRUuTj1
l4W9s0Ju47rxttoEPzhAgJzJLpeUYMRkw2r1RFvVyFPOuGq4JwFay4eK0luV1qCCMLwrADNjf+eV
OfRtSIxoIbia+Xkd8YCOgirvTLjp8LzHOR81aiAXKopod2/ql3HeZgAJ128IN5JXi3TmlwJL0IbB
4vz4UpMkmqrK3inELG7dX0xL7FzxUFalGL/AKFzTTzu8ztotQYt2tnEKvynv8MfH6BosSLjaJw7s
QKszQuFC/u/rNna0BtR2A7RlKZ6z99166RO6busd3ut7QIkds31w1zOAeyI0qCr0zogaeLqcH9jX
/nEBGOBzRAnmzBzNlpnm51tYsdP9DM2C75I3mmwIJqk1jc8ukTBlW2C8O3xmpxLIULZd5+yZHTLM
1F4g7FevWzqFmFIokFUsOdP70YP4WIUx7IQhVxqzxp9jyW45Av0mIM1xVluFECJXaAORrRI4snvW
vWA/N9qh0SfayG2PpscTrsv95OMFcztcd+e9q6YM9UzPXBzHnhsP08uJMMuARBJjI0Xe44+cUrZy
/Q+kcbo3vABp9XibBu/XmFTpimv/D42N02E4vJWMsATbeHDCt2QlBRaQITUt/RtdKkNpmqwDus82
NoeP2aEfnx3FjjQ+St7FKyLW9oSVeQonpMaMkWh+mDE6gjo0yk2vpyfn/eLTr/iR2NNVDkpUtF1L
sPEqA9U9h3b6D5uP9H6mBoE7DcqSpdTGBRDxEZvoRL6AzvBudODN7ygrxuIMbM2VpCdRLDCub25T
r1EGWQ/Ad8g4TaImGsAbm7BWGXf8rPyiAuYPQHaoR2E/v1wNXJi7TC3pLU0rMiBBPzxb5OW2TqYc
mq6WZXTtB0F98b1Q13bEpwndtD6IN4nCutJX6F152mPe3ZxwSdC/qEMBRMtrtHi1/2lrsWx3JVna
d57vLuKrqg6sYXF784IcfMT7vwNyS9rXirkAZXeneKuP50mOnoKbf9T72L9rmJ+jf79XYW8ubnNV
AsgOmwGlMiIdUHbIe80RlxIw8WkqcL4FF8osIIPGmXebmE+TECFJxnfiQ7rf/Sa3iH82qVjL9+is
0U6TNQnlpnEAj8XrUsH7K8WyQxf5q1Wc0FzGTP2uONkfYJo8EcIG9qAOPl2MNMmo8Z6O86uf/2UF
cDiua/evnOkj3IE7qhTTQt99tpCSF8Bg3C+wC3kmQAWq09WqWb0a+AziBtpImAWy9/MtK/+iLZGt
Dv7Bainthpy+YALrdpvicWHPAFn2UYBqWpWCPZ8qh02BDM5UgXw4ZyQfZv2XCRWg3NXdzMS7ZMbg
Cv7jAKM0Ac/1tmRIJHeZOA0N51wsaWc/dyGxRKVfKwP47jRlecaCA3n1J4IuwjCYlHrnG4ksbVOz
SDBaIL3+8r6jTuG/Dc4wCgmQKZLEDbfdZArk4dlV0DBRcEWrVvYcyd7AAv2u66xoaLgzHv2d9YLX
lH7ts/Vj287vvLNm+NFlImYp8cnlsDOVuadb3zBumG757BbACoVXEQMoUOZJdXZWJT35afpoq98x
6PpJj+Z2B7Kfl38P163g7IyGO9Ab8GnoOIr7rVk3IL5D2lbnKWkE9sn0JElGSFjWSLoMhe7aFnW2
W7s5Sq8c15rz5tdN3Jzqx2h6mhqBAZrzfp54lc8u2vOZf38J/YfrNH/n6HVPwZY6/7ez3z1H4st9
2SQ/4zW5v1fKFCZsosxRkK1YEP/3pPqHuOjgZNqQeWf9ta6FuOMGeWTopQooWRnqqa1LLSqvYjjW
JYWiowgwtLMt2uUPBHfHakh5eDXhX9hJ1UyvjrHfvAZxJPDy6NpcPi0ZD57xc0vzOXiQ3Q40g+ON
KHu18Xx8kQnHE8K+nsrwWUNz8x/g2pQWC77FFw43H0cJsZ68YhhqD94DJEiopLFqC3JLJniDrnHY
O74lMeB093KSvMh2xUQfHazURXtlZL7ExlEEQR1+4gc9xT7f3QypKUqcaMW/k4JXpeRuMHvXnt2W
eK9b/aneC7YUBVqgrMIwCuOCuJxtaLEl9EC+hBAggv8dlg5Cwo9gmI3zkVd0Gb+H6up+RhtG5SO7
d/6Y/i+VNY/1itCdRt4FruSy/9+8YJCJB633XJR1KNN8HTQ7Zj77w7FkoGxcrXQUfJl3wgf5KsqQ
jL13/002Z7ew1V3moXGdun8BEZeZUepwBJaFEn4utDsth1bbZhSBhDG70iLDQA6KG9BRz4Qto+vZ
jXJ1Hj31l2dshy4E4trqsaz4ZoT6qQ7wSUqsVGlUvy1DmtLhRoJjmPKMUOD4mRjvarT+IEhAPMxd
KuuZCUf71VYLw+qWSBA9gKD6KqiU9XRv8zgwAHOe46ow0wxkM2/fFQliwGn6TlM7/nNDH3w7mJJH
J4jY8elKPk6BoUYlXmj9/g38Nf3/AonZ7iI9RMW6GoH1gUlKKGSCCm8z8a0i6Y5M7onYcs3YYBVp
nVzzmwb45OLJ3bGMhntfJYWcYwOh2i0mK9Zf7J5zZvIXrb1IvNf//tv6Kc+h823ehfmo+sCiJSBG
/pJeDkdOKdZpX6hEz/ZfjZ/Uei5l1clbdd2ke81dC2/j0TM+64KKcUgoSfXw3kfr3i10jwQZ766A
3P/011QSSmfCA0XIndhEG31o2mBFiJtd1ZZ3sVoVYGfu9s245P1bWlvs7M37qj4U7aOGrtSuz0q5
sHdOydvjzRdO6QP4m7UYi+IzPFcwwsqCcOQNcXiaxmXR5pm2gx2ECl0+vMRvFXSMDQzg+l+FprAI
cnqjmw/yu3S2QcTkKIzaKkiMiQOscrf7JzU1K+6g0x6czNzNmB4eTpq01AfCzQhtfByGwormlyiu
N01VJFz61teYKNi7sWRuzyEFQk4SxCNV1XTKX+SBwrk6bIeIReZCZ8DXZaVm2pDfQGbmLlWMrVc5
1djYoZ1/3yWIChXAxIVMGmGliM1GHf1/M8AFCwV+k7wxqDhRwabmJ89fw7DYeJVUDsyvgcCAXeI1
EL1qSlTO+lg5GTaz2tI4vCwDz7L89o90pLsUVUjFx8Ff7HJoLkQWgxx0GVmYp5qHoJx8CCx3sEwG
5VMsBWGcteUU5fXc+jyvJbqRA0AD96OWK8nvWZBLlaMgccsgzZR1ttIwfOYJ8aukJmA7h6DBmhQ5
AbEyg30CEGHzE6fe80wzB9HYnwXc9SwKP+JfjTS1s8YyC+tJfQ8RSFmucRpqFxHlVjKZwcuDoT7H
ohBr71qKHAqY1Z0cL4Ef3b3D/R0YD5LFK8vNtiPlBOCyU3EstTSCVUqWe/mMim4reu7Rpg2UfUO5
asIL74FIA0k6jqwzRL5cKwFmiy1Mu9kPu7eRRUFFNnyR1PKDJ1UZPJZFzphABsJ1om5Z35XHdEWR
6nm8HqmGkLb58Nlxv+6GWYWbZkBqvZ7a+RkPRRD3EDwhpfFhzLrVHfvs3ulrANe0jH/Q9P4G2FmM
XE8M2bTCK2tgxmYtynT6sopFFl4BDO+katFMcvxnVYUeIomIL3eKlYyHfdCSPZ7YS5HE6K0UgjD8
6cq+MV8dFTcJnA7SE0Mt9XHx2fGKF8lfa8F5v6JSPlO8rs9taAGC9uUXqpLAJG74q0rF5TCcdt5o
I8X3ow0vCErvAZ2XxKSBHo++YO1ni9s0+fvjDQE+qB7c/nryPQlQDSP0MZrAmwhFwiyEw57+0PkG
cCzd2BxMfXkak7anvnMGSCXyW9ej8sFbyFwtMR1ZvcrENz0lDRI1zXxCvt1LG4KxC2nkon1pcF+h
oXn6syQslvUd6fNHa37+TG4OBdOZXNPj59VovNfOvHSkCockYAJheIH9e/ztNwID78/TsAuAJSnE
d7iMwlZeTEshSi2F/rkE0SRERjQvTtHGDuQM1T9cMyzqnavzMmbaYvXMxtj4otexoIUShhoqrpm7
cVX3Kn+aBz+yRZX+lGTOU6VHsxBacsRNzIm7SaN9r+SWjtYLv9dLXEEyWKA2093tvW0DOE2iTcYP
1Ijy5ja5vcX6xftJqZpgLSSKiKkOqmhWaQbuahN2fhcja8gWQfaXAQrbFGLkhajZqWRE3Gkr5Uxs
yAun2tjuoGukQMH2F83UmYcqVBQmfG5E6W7CSr29HRoBqMmnIkIAS2eMN9aj6qm1h30T0PysiV3I
MAmH0IN46iWpo/4lKvXzjPHa/86TAgOK+O8ZTgIU3ppvVwCI2uGjYGloy2Uby/KaETvwN+dorJOW
Mqu5ddOtTeyNTUPr+JUznsXpIAPW8hOrlA/O2ypUI49CTkRw9VR4wELkxSYObATmj75QtYO/9ayT
f7jneq1qu7Y0NDT1lPj2MScWZmryI+8+LW8uF+vm6KUPlvr1sP97lHEZFMwASfRaqiybl2e43SBI
SNLQSZZRGhstZXqM2gplBgydAGobYq0XwyiRaLbAXm4MP/BhPO08YLVqr+zlz8iQD9eAkUYWpiAV
hKS+T/AS4oGktckZWlxEfygC2xwFmI6fJgueGPFZ6zJikmMdS8tGdl+EVp00kHu/4G+XVG5EadEA
IUy2ahAzHl2Qyg6GK7v5NpT5pYWVJIDRjOBCpWVbVmj2lNG3FnS5JNpbN5zQNvNlZnrLc07PpKhF
CxPdMdFy3Y0tHCP9KdLVCsgSgQuy4WEwAaii2QWhkKFjDK3gTD1dMoGw0LM8w+gDDXBWoYDwhyG/
LBgN/J3ja7vGVrVVAsj4UgdkXkpf7ByNq7Z1sK+Ay7L8igY27x1A+giK0MMmjHS5SFgZM50EzhxQ
GffnXj0PpggTIQi9bNsmO29Zip5qfMA3E17AJ/bSVXn3YNyrZtbosrFmvSiX6qOIa8prKLiQrdfg
YB2DivC6aeYFGlYax6klhppbbqhYElKTU86F3YKJkef54Gtay2pKeR5OswhRSLXCf7q5fYtWmqWJ
hr3D7nmso9UP92PRCI7l/0Rz4Lr5ymtY7Y/HUOU9V6ojJqBPvgjUEM+FDT42bw8XrWF/ri5wUpIr
S11W9+ka9gMmYGSZElJhjhBa0BNP4nmAhOytcbTtG6jk5nFqbyCF+iWtHUnRz2Lzd3fs95Y9ZpUq
vbovEIwyDrS5jrrDSt+KyoOCj4SeDpARw9LPIVgKJFqCiV8JCpKSGKPvzBsKXri1+3+/hgaYN1zR
dvX/0+cxdFf+GgsShCpzdf3o1tJvdRaLX1//e7WkSuHVb4jqf7xmw23UUPvoCQHo7Dlfw9qt16jR
YnNqvE/9eyw27AacW7BJDA5VPk9u6jsGztDN6AwaxSsnC/zO8VIbEl8t/1DzgopvkQBnXixyvjZ+
TzXR1zMJuUiJFiKI/lDMAe437ic9zCJjChFHFfstkRQVjet8cGyVJhzju9MKJkdroiugK3W7kfUp
LwWkmFeTThcfishi/H3hE/77hjg3mVAVLbH1y2GH2TR4uebFiQBXOnW/hruFHXuPy1gcA/OZa0CN
ZkNcjcE1CDTLTuwsiVdWJiZPw4OsLnOYaUUBDBVcXNbd5A3yDzF7YH31LlVtb6q4erT/dRQLO9qC
GDEhvLtVLKiiv850CDCvo4+qR7JsWqIZQ9q9DSqPoKbMnfPSkWwHyEEAWglGCfWE+nMJDCrScTax
38RosRS2Rel9a2bIbKM2+rVcW4QR53ZWL3mHgCsjGwmcqeeSdsRL9UngF2OaV0V7f8fOYN86hiul
pZ2GjudW11UjS1XLZdrwkqSGzxlQ+y5Nt0at85g4mRTm6m5aMEodF7CzNp5hQ2MAzDhfjtDwLgfM
aeB54yzUrACawJhvdRzMH69waqZCNbqS0Moq+EUmfvTcKPfKL5K5MXSQoXcUvSK6XgjUpumIzFHy
knfO1ZJZ9kOAXMEgW0p7UkYEsQu5/HRguB0QYO4lvg2xWDcRRgTAn6HLf/VjQ0OpSgMgY8ZEghXF
gMfViyUrRJ0ga0f6VvmpZslJOnMXf1m+//fLKrKBTLS0NvVIJkY6Ytr2tSa/TjVbClZuARQzXzXZ
DPpWRPzRhbsokA5DtA3iTyj2hhlPgRlwiD+o0CqbRmzUGQBre6qGr4KedIwttDGZlstRrC37K3yR
4EDuuWmySi7dcA6yzk+5eM9maKXz+9o49yfJf7nCct4VfguaNBa7kA5Yza4m8OJ9T/sLtlbFwspC
djcX1UYgu15in9BV6KCarMn9rNPGgrk4UTuTYokmJAHF1SGScHJOHPeLrBPcuz1eDTnzWSdU6Mns
Xds8gQhmNbKTYKt/78SxtTo+DIL8LPJFWX81ePZOZ+d24dayOMOecZum0g3It391tjPsr5YC1bP9
AdDkoGiPXtREgTMFbI0tDxjVosLllbaHHrRoV7a6mdlZmmuq+kFkOIheWLd27sl2jDjFUIQxMx+5
6Mv1JSWdYhzOa9sW0VY1sluAJ5sxj6P/vHwjeFTlxebcmzMzkBB0hh4AaGkn3NDRcw+XR8kq0nDy
77tLmcXiatzmNDPRLnBqKmIIAVnd4s5bH/QODXGqObmrgfNyniSYilAKDEtnK4sFKsk8QlSnByHZ
hqtTToZJAluyAJNhJa6qgCE9gQdbd8nwtC43RwptIikA+6Rz17nTUXgF8vHyHI2NlXuJJwXrJjFx
AGfSdtX1gDwOa2HU1ryOwEQHDixe4pA3KJMxPzet5XannhCLA/zr6dANXHUUJKRWmyi9JCXcTwUH
URtib3gBDmVKe7r46pb2zBcWpxhDiprM4MkVqKKl1vOGAc3VihpvUQIYJkSjuZQAODQuiZfc5oFa
HZp38e6bM3xUYUNCNn0KSXYhiEzdOEc0rDc8gI7MG150bvJC0/rsvQgeL7w/WmfO8NYMBDhsarTu
5ctCnduBAxOzxw3MRrm1GDLxsROUo2LzzHNdLPHQXGyHRSKhhJEvHclt1twB2HELZZeXOJe6Qq01
u5nysHYrgxnm5do4t/w9ZBmjr5QKM8uAQaqG9utDEqJv0WIU6fWsdTzbn9i1fP0t1cLR3FGiK+Nx
xT8+LCWlnAttW+/6Ka30bO3WD7CioJI+I4Lj6Zla+qicQRYXgd63b5YIJwtQduGYfiywLKBYho3w
NeZKMLr1S0NwixCubYZSXGJo5S7/X658CAcxB28TcrIOa24eUmsS+I8NfOcRNIY1XdVZ2hkAZsvI
rUZ4S/DHb0UaKeVgtOuvqAWkHPr5emw5ZODOgBxPUXHx7h0esG9+fHfP+YrTsNazYs5Sbf71AgG4
xPSrH3KVdxqEmvuQiF2FI/+Bmx/u5HMXf9liu5923LVp1AYf7D80sbljpGBQtccTSA+eMjjnGyxy
KNhjSit3NKarQT7KSkRaaOy0YFjXBuFrcoIJlx1LO8YCDEu9CawK42LEg6IpZd17+V22+6SbAQ1T
6Shu/M+JZCCQVu6Cl/exwUIeXwPQUDlPYLB9atQAlBw7j1zCjldk83Kh/zdve93xQOBFGAJr+0Pm
/1ljFAnP6yn8BCqOKOsc3F+ldlaAmHShKxenMr63rcUDdutbTItalPRMweVIgBjKWJgA8P23fRc1
0Vv59XDBt1/0LxBZ9VxjyVt/wn4M9TXMOlbA1H9t15X6QXvCVJeu7m5m2E/+gd0RAMN0CuGXxfi5
c5yOteqx3YrrsLzCQ0YJniGCFLFjAnkC84Qo58Z/37TSm1yWSoFMwovr26JrN6bX5ox+ukWuEWcA
EoAnnfI3IduhCtthuixRkkZUDOy94EN1CfMWHbkltZfELb7AwLBIETfvGIlV5b4KilGC8CWRxi/P
I3x7Lu6PKgly8DK94nbhZsK9vveSl13Gu3Ox87NHKzF6BidWVfsydWk9UA7lkIMNqRaLSzCveSCC
jhtzi5qTRWdZNhFoGRpppJcmkpA9Kd/aNQkaXVbJHqyX5Z69UtdfexI9TEyGBl6C0aSJgKz2lbQJ
cH5J/Npo529861BePBNqINRDB+cbiFYGiBXxQEY45Gm8LOMeVQeRNV1fcdbdNrg7EoRz8vE82zmH
0VULRf+avpIwG/QpEmjs5y0jL1s06mumqWwpGuYPXkbTE8En+J3RCSndP0J5b/KvqaqLNpDa1jkm
yBix8Ntfxb01IkxQhZsYNYs1Zfwc7l1alhwd4mZlzCOGJTy73f/CeHcn3R6+XDS7dNFIw4dzOBDp
6cZvZN5Cjkh9hgNMXAYRAeEwC1DmhMnybwWeKEb36/klu1HWHlZLTcYBah1RlFCPIiJOlmLs4TzU
1Kt0xdt6IO46cwTtP/Xm7guFEleCdfZyST+ZMD0oOEXL/dZn8rNXzPWuO9mTlXWQkR/h5fwRxmsY
kOukK7QUNKgQ7I4oZRRQOICAGAqhjOGPn3fuWYrjl5cI7Jw2edLBbThkzUeYJihe1DPi+QNMbbYV
Zn6JPwAQXGpE682+huf1RT5VLY17TcN5J6Lmam7mip1AKjgVjiGVuuGwfu56hBhaQhmbE+p0pgf3
Ul621QSt3P5MpbVVhzb2JqepeukWZLvk+5mUNNfHaZxiWPIrOKxere/c2J3BOYgB0HIbBfSYAN9q
GeIlK3T8A+9nGFChFZpVaEoPJKbcmH5hJRmD8zGETbMPAyxPGYuNsiaoGRxvWsFPrUoCCHbOHsfd
PITS0eoHUDb0ZNjghT6y4fw3nK1piBlJXlgTvjx3bIKvKmy0cKLtwbX3Mtr9u58adYtE+Lp+m7N9
EQ365Ju6mKKvTdsAyN2JGH/rU0PHHCmNB4H+BjKAG7FEwNcBU/fY5wctRZ8KAeqyL/XVJlcZPJLI
vkFyV14QGX4AQZp1ibqa0bais2oLpOjYIGCL11qWmlzc/BV2/uYnjHuR4whNH32mE6zUIwK2kis3
NUqYWb5Freaf1w3/Fk1T3k8pCtYm4BRBAVdTjeBvAmqDMohN1v+Rglz3ObC1A9fQDQAlurl7Te+e
FQD4ieYim/8M3tzMEirJBZuqe2NHQ/B/D7ymRtjopRQEDH5XudNWk8A17KLflmBoPCOt/IHsmcib
EBlyn3fmGoLc/n9CovTg39TccMTtA4Bi4s9gRiakd5TYSOkePI35jirKp1SUKio665mt3bxB58LL
JuN4IW3bDAPzfqOmwuR0YjtajCBIbyM9NJdIsB3bvXCZoU5ERQHSpzj4KQeU0J9FYKwhwxSP9ABj
Lt/DFdB9ppuIPCEXsieNwFCuS+sMvfXQfPtar6bUEzMQwd/G75mJq9qODBi/z7kOWB0dlAQwUzs8
Z/QGBPvlJEqPOIVDB2E4GfL1Aa0Tyimazp5jeEhh3Ozia0b7+Pk2LnL9K4Gn1QLZoUpO6PpX+xie
Hfe1jZneBh4tWpKcT3R2W51PkkA1sSpC5o06t7c8L2LDuf02XPvtsgbM2ObgGRxkY3qVzR+aAcJN
XbVxH0REiDTFbLhAt3kITh9D9EuWvDQFpFmkgHXknZgTLK1PRCgR9ItXDfqLk0Q5nOPVaCqYInd6
zt2WM2DTC9+u0Tsqbek90gTnB7VUI9VuiBu29Fm+TpnbwHqbXkGPli/cAdqZ8exgdaNoZsQeTOby
uNwwLo98zjNLAoy+j9yhIRL4NKCntjOCg7WTQa/UFDTek6JcFH52HDV2k0ubRV7unQAz0sL0ipNb
DUUS+5SDTyTBIl059cgCMHIee70K0f8QcJrC5pyW+dzY2eIeFYPpP2v1QRA7Qd2cHOU9vwCbwAr4
Bf2vbuZ+2xCPmlmBAN1f5/8bBnUel82NhXpl4N7Mdu39g4nUFtY2acfjQNmv2F6BTW5BSW79pc86
h3YkxVFqsRHVMKLOK/aKwB/UgpR/lPy4iSVRFUTFH4UQQiXFBUz09OUVugU/DnTmi5E0bKrGNxtC
sfD7qIW541/D8I9qZdrC3hQfTOKOQUI/11IKfPe2YXUiWpbpT4KKamwzNW9tvt9a//E4QxnpXAHf
wfte6ft/TjXZjXvVNP3cr2Iq4XGBpesBp3/rP4fSjRCF6KpStzyhTG6wv+amZ2EPEPOmVlP3JRGS
hvsqH8/DRly6Zt5mRIKj7xZj+HN9xIZmo5378mmqmM6cw2U7oO+Dwou3jpobDh6RBod3dkAmztfx
hyp1RpJ4+0BoRaZ2u+b3NLL1N7TzhrmD3FhKFNk3/Yf8GrCKxgCTH+k1MXdL/xHmNckgUEO1O8AC
EJEChHrvDqvjGTWrEI/DKJI6tPPZVsA94RuCpywyLgNo8uShPa03/LLINuWIcLp6nRImeFsUOeZH
VfnQ3Momq3IHvk/HaFG2vfKzFXdpMg4Q4X7kbxFxphaXIm4V9/rE7MfY0+To8hR4iONvA9iiYCgc
a4g5Y0ny1sLYqti7HhPOCY8QTsjHRv6QDDTXQwpEjRP6SyctCu+y5lQUYdtNOvJySj4nzrphnWrl
qSvPtQEL6nYFEwIJCd1KUlSivNEwzi+Qy9wPGNnSKCN62n8GtXClmGJev5E/SummIzf1r3bpI6Az
bztzPKSJmz1gvIvSnaag2XVyNWXbQib6YpUVAPx3dNxWyu0bxSBCP4HpvBhAOI7qWKzDKiMi5l6w
JNHflGk0+zc13BgL7X6EYDKwuPtJ4SEdtD6ju67eYATKrKECeRlVOCxuUs/77CeufO30cFq5JItq
w/2msP4vuVzX2X08QpeEbLE69nUHGHl+jUslduZ8pj9ngSuKdMzyEn7N3kDsRLptZ5TqY3Hqr4Ju
kKLPVxVrRtZx6CN+7IEdkW7SSjq55Gaz3GlvOP+VFmJusCHQTfWpRLLdx6oyZ3h2YeBmBeQRbyPU
8708qyvnJJlhV1IDDzcWviDBkhaZBsYmoxmwU+Dke9dTL2V/VmZg0YnngvovIEYWVUyhq8CeXEiV
BG4akC40J4wK/3uucS8PruCQqEjebCLV1CUJ2L5ABB+NRBMYUBsp5z9uZ4t4JL0Qb8mXYq0cZ7Wk
H1t8SlKPTxFseKCuGfZ6Yj8bHiN94sZ4D2I9YbioIlq0ejVHWrzTRy65gvJ04dv0zdKwyI2d546p
WwFpX7lXsU//wyZ7aSvkhYfY4zf6UdfymkSpy20nquVTxjoUsJ/4d7qhWgO1KIYgBiQrvISwvJr+
4VOYWQpE/urql62oFXuqtbhWZEhMPWAxmRAWK2htbU9GH1NGKFwTNXiEPkffaeCS2EXtQ8dqxhM8
HPeQGF1pn6x4C1TbOMld9J/dWl73uQ+mIhGXWq1pmBWbe4+v2jngucvj4lYZDw6sRxwvtQ0VOn8+
hpROEJHQjc283BjcbpUQC9cWW4b3nzD+ynavfSZkFEf3bErZjcBxxTiVdovG/l7r4rySNHckG6fV
IB/gmDsUXR9XqgWFxjCAJ0sLvdlF69w+FUxghhU2+vKkDy51caU//LAomkemelZNN0xZE/stpmX8
qehzfU6lLkmPpKG+x4aD9mSM5Z1LFdkCYBIxcc+UKQkjgYYRyauyzOeuLPwMEkC9H3YRvts9ov+0
8/1ZEhIyIsTmDTOELyYoawYVtT50CQmEHmZanoTkXOBGLT5f7BZXr8y6jumb+phrOk7quzOliAk1
G7LxpYXzXnOkjwTqqY+1tE7kCLNuSeYGcXzQ8MPa/hXAyN2rndWSkMt22ziVtVpw0aqlp5yQRncr
w4Q7gooapRTAXAtbN5R5nXgb+SPq3nmNSvQVdJB+gEUCmeCIbM8oWvk/rSWMALzZ2Im1+fNFQM/6
NMjuE3ijnJ7SMWwUjN3qnZEKNoQbeknmGvttLGdjY68nzZsh/bqXakkyukl0bK93bPqiOpVs+Gl6
aL6EyGXH5n4zLJLBv79Zfpbk2AGK/xQznsSyzFpFLeyJiL8FBIE/aWQTvfvgdV7cpW5mTn3aMWti
6Xgdck001iBhPM+v75ZDdT2wNpVI1V0ZbP1YOG8ya9PRUUOuUuzBPbycsz1B6iO5kvj1OE1Hmzku
BCsNSxic1lvWvc8PNg0bkfq3iAFzF9P3VgZXKUNS3pBPgELTMxLfKbZfNRUL0snZx5bIZJHKe+Ae
GS8xIkFDdlzdH/efgK31o0n0e+VPFnFRHVR6AROU33+4YO6MS18R4inFK+ms/i2ASjYl98JJHbLM
nzcX2XCs81U/AqZMmbS91Crs/pEPAoW+1s/tIJZRqkisX+GQB/LryI1eCfIJimjyuoeSbwtt5cXS
YU1QkioO0Xwjs64/6+RaJpCK8OtXcizEPVLdFnB8tcxPAn1Nw0knNEN2UeUHV3sB4JDzvLNTrCF4
ac6B1IZZjcC6rFmID5ZCFj1qL1FXbG0QWBkuuHYquxpRIww6S5OO7Cg5TmqDVR0eudWjlpu58G6c
x3FW8pVUvfpXLRqTgxQAsypkkB0zOE06q53KMaykZOnvu8OioUNDCq+4DgLrYmN9fcIv7ivdswve
k8kGmMqmZd0RXxomb5g2bsOP6FtVl5qLRuxRTyoJGtRpZqhoqECKqfZnEmLSOx21cQQahqfasDhp
QO6VBqkv58EdJQsNNF3B95GhgY27V/z4kNBldqXFnZFfxdJMmgQBjMt1oewG1wUgQpcCR/H1dRlW
KrRvRZZZ4CjkEOPpiCF7M5vG63aAlJPyeyBeTiM2Og2wAv/3WnfsWCN9i9d+mmBWfNEwsX6fwx9L
MBewNT7dSLcUm2MJgykfqC/MCpxTAmHvEVDDnoDDupSOCy3EdhKTAxnG+1MJTOAby8I0/VeefT2k
rFY+rfOqgWxBLHL0alBGYmmbZubOlmlo0mW9kqxeXPFG6zhAY08LDzvubQBJQodDwYRxCLPFYHPC
JQpHwdBINRaX7rOneWVl24ZmJeCeSBkM/Ef5AQDLMC107N+UG57uREHPvxxCCOq9ZG4U9lg+u0Ds
oGM1OYTYxiePzCxwmbBjXdOVa0tfoBT1jcEjWqvc08Lcp3UzetaVR7HbZ/l+Tan62pm9SpPdV8FX
NXmF8eXDr3OM0azeBXrZ/jFyb8cy1eHVVHEu4+kLjThgLh3BEPZs6P5eCgLThSf669YQDGg9fcDn
LfbJjHanAfjEo9cnVc1jfNaHS0Bc8rRkB1yrTxBQ+FbPfX+Vmez70C3mL7gVwuWJeYGSlS0GaM4z
1TO80+BRE1mQ3L/7n5J4ROfx/9cXfpvdcO9Xrk2QB4Q1J2+tR/28EbvaKIwVF2zP+X/VzyfWSBA6
xStBDTbkbZAmXO5y5tSnZ2kKGFmgsXNZfBNNNFCgTyGVX/GgWNUysasHeLK66NDg7gU7Hwaz5khB
cXMklreRXmUL/Dm7BurtNAeGNmSaXm3bDHwdjrUHU2Vjbu/ZSQixufBBUWN4CU5MmRJe1raDxsT3
BBdGikkLQHakIcZau2dlBjiuD9eyEbPC2Qgg3Q7aS4PpeOw23+e5utL4FztKMDtlhi90E25un0Lg
6QCQRHs9Pot6YQ2vuQalX8eZnrau5vgjZVIelf66pt7aHqXcP5HjmDEKYINavq+ky6/Kb0nvfy6J
fU7AI6gM0rfaJ6dpQ6noX4IsdMYNA0f/gGR7Pkg/B3URHM6h7oB0Sadx3J2NmWx6zstv7BiqnXHT
KeBtrDfL2THYcWTZ8iO/B2ykfEuNDds23gsV84+V0iVFM2H6/XA4hnx7GJ843ZxhCyJ5sUjvlcvl
I6OG6ZgV5gIxSGyfyxyIyLxcx6+4bsFO7zPchDwyAXFQfVG2dtoRORAxr2fI1dH+j0uwPuQKXSbw
y/tMcXXK8UD3KSofpCHnFBInZQzV+2xLy8fWuv2xoM/FvrIYIKrUzJijppDh8NLSFWqabn6bUAOe
iwbWYej0YXJBmhVyx6XcApkV4f5phcOu+LkULH4OK96lCxsf0/SdQ4x0xlpG9vxUfMecEVbPdrUO
NBuW7Up+BDHnVZDUgcvj2xzC8zH5q7uRu/cPpOLQ65tUZJryZNBpMQs8t5sdC8o/rfNUDRCV6mNE
vEU2pP3ycN66QbcgYxk6WP2R3Z6JJV/BtmcEP7l4SLuRSUDVWzV8MjzZPY0ev9/zTzI3eHnzMBWu
ktjeBwiOhu48cWRsj9C4Z/5xXVfXICA83REeWDZK/fOCknpZLzZbunfrxLxk8Dh37s8u6Doxzlaj
JNkmTdwixvaBly5ZPPD8KqDpDgpP9RDpPu0XcY1YShYBxb9iiIDNnhUltMtpm7TPdtoARxE3mdML
KQLcCfgdns0Xp5/tlgH/08aOnRhpQIIIMK/Ukv7Ro/s1waZ20r5WM7qfmAaLGMbZmB5o6M4TENW6
vdpC7crXOkqkmDzK1dv89mx4E9S/Czdq9XRUOe2CaMjSjTpQxEWQrlDXxBeShOhHSlNYF5GEiaS7
fhARgF7iYBkCbcQAlG9QqVXqjuc34a5eeiynvqwtvDSXyRHho8p0uNbu8/Mnb9oRXheHBAtgFYic
6d8eggZS9ad0uReyuohF467lhNHR4WQvLTQ3peo79twDhaNluA0WAdJnTIsBG715tnjqgH6P6OcJ
QET8EdBqg9jCJnXjM3i+OKelEh4ftO+xiB7uQJLKPHgEyPKIQEePr4mLW5T06zYVMsZjTwlkqgxL
JLZONqJFe7wa7Lz7FfctqffstCGeYOSesEOhp9u7WM09+MXcn4zka1lyoqeixqlDGk+Ojrd4TUom
Hp/7d4oAJvynYcp8bIYCBnr+EctR/STjzVTR7uKEhG1sON42AwyQo+1GnGlZ1AbfW9S6MNepgP7i
t1VIVmiiWO5P4CJDzT46xLxF+Agcdr0uQ2lXIpmugfZCbEx+WjYR16c4xO42en1AY163VPfPSpzQ
7FIsGMsryotSMy8UqaE7HDGgyNuV+8XIT5HKRPq6PkX+ywVfC7oejZ8V/b7fCyHyyagNQtATge3f
a/M+0WG6a6rXlfbJFvX+t73zSAjdIIBmC0f6rCJkkK1Jpuhqq/5DSyBwAjoLuOy3M4yLUKTi6Ld9
0aeuTpKPrbsOYgWLm4jd/nzUwl0fvP3FP+TnEMAYvcNrpQJd4HnyBidxR3QlRJzbty7+9zBHffAr
SQ6OtNPCUCHfx8OhbiDULaQ5vZOiMF1cDwDC5seRHziFRIDPx85DxYodFm9SO3tS3dWnFQn17FFf
ZTnbuz78f73taNaDVUjAi2tkQ1lQBBL6k+NqGboeQokM83rR0QM5onn0PIbJxFPY7eu+lgEEJSnb
m8S1nm7S09lMCTw3xnNDyQk2C9e56U2uX7qREzFX49yGUEn2medkgucJ17J5LgX5aEhZHWLzKhIw
caZL1dmRBTgejw0zGuFQWhe1ZOa9E1TwLi/5rZxmFUI9LtGcflw/7Chyg7EKq3A5M4HhzforrEsL
Sp/DRIwqj09y9VKJKeoH3DQi6Am9SFBRZWb3g1yRlAiy/kAfFFMXAnNw8R2qveQO/APRVTdgX8f5
S3BH0F8m4QSGNrVS391O1cmtYHmwb9zmA1NTSuAjnY5HfjWVo01U0zuMas1VuMmrGzr8fSaTM1bR
xvO1U1OdYANgstMo/hHBglWTYkI3FQI2jK7VbLhdpl4t6Z5WTuXewJJwkxS6AenY7WolH01bH31k
hZ0WSuSo1CO2sb9+lHl0bn4iEU/bs3We+poKL0nXBSZrWTq6f1ykcrJELBzdz5FCsICvQbePYPGQ
kALo1wngPQI9fbIjPKAYeIvbgQmNAPjSTCssPRO6YZqyfnq7iC5uiUdcKXxm6DeeTJPoM7vreX8y
2mzmiOzLUcAKp9Pba3ssHFoPyGRZkM4LLHVSx9vlZ2PMWhhZ0MVoF0rWwLt67xyiZNPktWDd8P3b
Gqh3RRrYvr7pr0HYHuXR/pUw46gbFiYQ5JVWE81WYhfdDX9Tp0dy6FXoVcu2ZYdKH3F4oK9mVwER
x90SvzABj2SkxnZMuNX8nx/tJQkKThcS2s/o9mO6ReYM2JETv/fATiaSzPW1SVdbs7uAIpX7637Q
+8//4bZms31Ofmb5BKNuRILQ+ID7kayzmoj9fW8Sv2pY18wyaFNN1FLfu2UfKV2S66L27rp9/a+c
DHZ8fyFlg5I7ttoPqeSzbCLB2msJdwiAuwnHkqRUu/po47q3xV2U9ms1DM0jVY5VDBZU8olq3YB/
9BDXDkI+XSVDWNd6Q1/wcivYz48Fh3CO1od+aCe5qi/kAGuAWoNambfU79Qkw159LOy009+YAt1u
sucbrL5eL6nR9HxU6emkSBMeIu177BbXLBsaaNpBV5UvQrY6jOLB8JH0csu6bS3dLk+v2BauM5Zw
Bj7tdXZ7Td9xDDf+Hc30UioPflmM/eejVkjYxNN3Yow4Lu8UNRwesniXIP+C2d3eTSnzOWrzTNL3
zAzIrmv57JufEj9e5x5g0mTVPzZAe3V3NniN8cdzYiNvI86Tl81bvLAo+7Vf1avSuI9mUmDasBbJ
5SNbDEd7oqar7kouRMxHvvsuT/0xzEPbyATkU2l34aRBXBFMUwLSUM3HckUCTjo4AyiaCIXSXjZ9
/f7HOGUqhZ2sXdEpVQV7L67CIVoZSkIJoRuIeIDB5vc3R3XalSaFBIPk+XFNHq7rp5BZ6uJTc/Vs
XNsLlPy0xeoGgvGRkHjL8d2X7RMwHL6ziBNJUtX/hJLwJJoitCdRpD+THWnZyzusutIA6nyhxU1O
DUxNH7mJPUg4M8+pdrUO0IX8eh9II776yMA0apWrLvqo9KX7ELgdug0EycTYVz4w3IO8Ea/P8+00
bl8ebAnPDs7jkT5m/VxswH58Diukj3EntiTSv3VJTZJiN6pk56HdXm6/qo3cw7PlXp7LkoHoqb8P
Rt56Cjc57mIHqTEnFlHmntsgueQ6oVnRt2zlelURHc8Yb9nuJGlwoEdFRsC+PgzNCVADk1V0wIOJ
MOrBWG0WFkmJef5sj1Viqs3SvD5HTCFJBUXeSYtgcweeECoPIrPPFTQ7/zvORGlp+kJezNsW/vx6
plyW28h0b2ZROwW8gGrV5yESq7EyIze+En2rtFqT7CAAbzEAJld+BGDZEcezGLxDxWZeS7pI9T2x
P1B9gnoJC6Z6FvFlcpP6PHEPacaYmHyTAANUy0iksubDmqLOoJaFNIW6orByFD2Bs6S1KysyGj+V
Zm/p2D4dFyeODcXmNWglQVYB8Q+nCuwD8PMTODHDgrgW/97N6rXdpSEQr0g8/svcghsDZAW3Thal
rVySOnxsoHgqHOdcRyflF0+YYGjNEXMYrrSIW3OY2hJ8coMeZwMqoQ3RBOBJkf+hbpJrfwYy1eN3
ijqxciaEwuUDTK8NLj75oxZQfWyXegt2XmeEbiKBfQ4QdboYsEJ9Tk2Hrat2rNAvSNpGA3x+zdZG
eJ7cROesjRlHQyBLw/LsyZmJOtLCHBH7EB6EFB3Vafbfp8U1fhXRQ9Q59cK65GbPGZAeqZ/DEqtR
EdJ1DzT30foKw1W8VHPLQL3YdQvG14QR9zavP7f8UGQJt/J2LYeHCy1AQMDgFXImEWopQP+EFs5C
s3ChoAdJWPPm8Mu5gHt7S0oYF/AN8WhujVMwJDrvji6tB4l7JmEaHbZ/uImSSyfJP8X4y9Qm1zIW
RJefZU3udm50ZUr43nUw8Johv+fHJGdV67p3dppDnWzpk2D1Rxjr92yNBzlCFNjyiGUANeO7fs1o
OB7gQvUJjNIj6H2+u9nfFhjsIa+HwfLKdAHs1V/kzqlDVybKJlX6GmJvGTA+iXDFHru18F2qtXF4
pMkgPdldF53Cns69DUmjupz01TZDh7NpZFDaTG9VlHtCMdLht7mB6j39be1/agXPFMcHkwYZQR/w
fLzvZ4t8PhrgJrqv45y3r2har3+Q8mh/ZTc2kIbmOIHAp5JMin7lSdtbGtRjt9Y7714TQgU30adF
q3fVySRkMap8Vxe/V6e3uBb3QJ18ywmgOK9ikFbeOxoA4lCKzz6vVanU3Hj8B2XA2A5th57G8JAR
9fNXMC1Ut2yQnQ9+0fTF/r3tSf14v8R5+fq3IlYqt9y6EI+lrvQv3C7BCPWcXzKMQdh4MkHloL8B
UUCPpRe9uybJGYam/OeVt4PK64TWIBX38he58U2O5lKVXUScWqXzQ4ba9uKcQBxQO2hSo7nUk3lj
NK7nK0+Lvfvb4Dbbzvg+K6Wce59wHYLb+Bae3q/S+11XsuREAFjUFT12nHFstG481UqFX7APsnW6
s7NDkg76941kMwfP/XM4OxKG6o0m1Fegc9Uzo8wuLIDPWO2DRyyroqY4gsaaNqD2bU2KoXVmGlJj
CQPCcTaxt+K+MAW6f8nuDqtwBm4ccHEiGrIRywbNpkZyirdQ0NSuI/+LRfP42oF9PNvS9JMa4ztn
oYEoXfWYwsgSC9Iepn7mpuNXfjv0JqN7bRw1zeeC2VrsIiIUNRHsd4xtAHnCEAMGlH0ZKATbhmgh
TD2m7idVVOfyMI/41m8Ya0Q+AwZD9s1FIiMda3Xj5l1DM12qlAb3oNvuaBRovcRgxTPzE4AtabQy
F6TPLfGhhLJodiShORgSt9iM2In68INbLRT5DAuvX6sRsXg/fyKuWEiaAm5F0BwOrtdcA1am7mpI
CXNvlDU6EBoQD3GVQSsj8sGynhD3Mm9WAkFjHlasjNVYWE7s6X87WXvSDYxYxjbmIii4UbjRjVsj
tMiXyz2ZRPmPlZOn8jZ8EV45nH5WBBBKgcWAFAKDr841h+oKu0+ITGCjUkAKdDzNcUNFE6MZhBdc
FUpfRLhQCigBSpFBQHQQ2euRhjSXTx81oCt/422zvTdScAKxmHt/Sh8N9Vg/ADCUPAJkz8B/5fuI
EZNSigK6cvJ567FkujlmAhtYRBs9zWidEFwMLuDO6mmANsYJdeoDHv+VRNwKZDCT0DNF8xZG3HvT
htm6AnNKPDgKl/I+eQEHPUF3S+nUe+b4+RKVyM9pZ1J/QC8qKzcji/AEiickGAuHBaAOuP5nXj+T
bOWG1PK+SkOhGPBvof9uP8rG8LTLNNasMFoKHC8YrEWqCc1l38aWwjyoboFBjzoL+Irw9Zh63cY0
lbnzNHSkDd2GnkawC3g+kFsFjYK1NI1L+6LLsI9JugNk5+BgMb7caoDmB5Rbprj268Bn7ecqhqK6
0nXVG/rwF+1LxsLyAvMUZLmWOyU8UQ+IEMRE4Bkm5ZGAQfgA41TfVxz6JIsFCd1XGij35lbZI6mX
QEK2hTdIYuL0n6MIk9BLkaNOUiVPRmZFzsHtA96CfRQzXFvutEQ8GhlGRgIESgftVAxg/1iiDhx4
KhNik1aSAoAwNUL5FSY4ip8IIu7uD9pI8D3S13IoEi6s3wnl30Akb+1/ZT4xnQlqckyPnuWGRIvR
OYyAFXeNZoEeIbHvvTtbc/RmHYTCjKkCAZypYOStWjagMkluY0fKEdf1CPYrDA8GwPelbJ/JKAsB
Tcz+FBMov0MF/0iePDQGFkjsi7K3w2jyPGp5kfkRjB2Ym7aF/a8NWIpqa7qXj183B55IugQK6F7N
texCFLTdZ2JmRGtFKRvOYzZtE8rWdglSx5DrXIvtdeRUSmsGeKMJr3csMxZpnJgA8QB4mdRuTiwu
PGw9XifF6QuC59Vy7BwsNGJy8bI84FSY0iEi7eaYelfEy/hva/6eKVTIiVptgdBslid21atBE/VH
RMNGIeM99izIu3Q7vnO0zKiev/YchtfR8hTBX8XIuKwFp8ESFJQIX2t0fxIYGXuVev/n6Nrei4db
us9i/toQFhvfZ+Yx6J8qFJMRoNFWQqWh8Dl5ojV130kExxoNu60qKDf9fWJuDBLbpLPJ5ZKpR8iJ
+MBvHv0uc06TPqUKzS/FuJ29ZEvO91jAWpMV8C0BfD2So+rgazHucsogQ+IbGI1gkPUVAB0U4Nto
rKW+BWr5uQqAGYyRHxTUSMYrVzKdjmIbIvgc+yvNac4jjS7YqsW9J3d+jTeiiZrk89XVDF3j55un
5FIn4GnSRRCiRJkAunt0j8YSAT6cB3xEqFfFfVgFqv9H56BQsZhrVzviAyfkj8pkbxvTDUfXTU0q
y76nC59nzCxv2T/c9YNgnXy0+81jHZH7uMv1EoDsMEGZnfw46J26FVR0V6/lStbsszawMC9YXy/o
0sQ6GtLvJAGrEAmc1wE14Y+i1nrWZMGLb56rHSKcsaGZfN4faFrXEQqoERECKhcXw888E/cjeSqR
XIry+83KxNxdDke5AXvbt3l9AmMt81KqgVUxuzS9C1MzXxPXHbMJ/12eUGPXbQwsNPjAVmAB06ki
IzfKfkBiiOIw5N2SbobcZf4+ZkqvcX/f3AA5xIbWWJAC62Wpd82Mi154jcrjnQhnFHzjXdrHOFen
Tc+u7hhjmta9VP5pJLEFot5hv9QJBAZeCVrWDEfw3QlA7E1uIk3jI0JuaizCvkiLgArW6WYOBrbX
///EG+uKRBnCAhsyA6qYWL1mhicImodBxTjQc5xBEyHAx6V1yyBesrafZZNVtiplR3nrFihgI45h
n8RmWxYjDB761HtcJTyoEN2xJDhabomj47Gb6qEaTPZK3Vzrf4bAGyGpv3BsJl/UrVj5V8d5Ny2Q
qAhAPoz86nryOcUW+ldogbk3ic1oqPkMTJxtUO7nQmnnvgUYAOra07RhRfP4gqHalWSisWWFUzci
vEtlotLSvtQfGWTMpoa0kxN+Y+U9uVHkjJ1PTddPm07t7S5jkCTvH9muM6J5cqwlX4tnnc/pUs4o
dU8+vky2nYBaPSg27LtYAQhNbSao1PCnOK7Q72jpbATGDR3C1TmmGHGxr8EFX8tfBO0qPg2gyInC
vpGw2vh7dUUCFPSApBL6w89oCwanbXRYB1afdyO7Yx0Yox2rxQLoc+mFMRQzyUmiNnvPcRunF3OE
ok0j0jkmm6SaBZdkZWpR4P0mL0Sjsl1EcR7UQeq0zdva9EhXE2okYR/rBMU7W1jHrRY/T73nrpNu
d8xf3cmR6cFfZxweYAgohDq6WUgVy6rc2SfFfhZUCa3aa5/YTeG1AiATr3Un1/X4ru0WVKR5/hB2
7fBli+s3rHbTwSJgLDqQPldreRGTuBp96iLjXueALkcesd1C4rZz/7SlacdYFULuc7pd5m3XuxBm
rZaMR/ZN2l1mPAFyKf2RPXWuVmJe1Cm1qgZyl/ELqB3p9r5MBupMqZUy99+Pgp85Lb+vQH6CfVvo
iqllGGlcsl9ocCCjlyH3rxstlPddxhJdOhUz2+e8E/Dha7jp1iRrZQdbOQGQG/bGkKYweutukQGV
eolLshIQa+8ZCF2zwj6E23ZpasWWVQfDmBwqfUJLlN/5IcPUMW8dENr0hvNDs9miiNvHpVUN75fu
3ZjgHV6IAICQlPk5e9Jb/lpmw2eBzlHKhD/f+JdXJxIg0U8BLiKGTPsQaxyE36zucYG8D8kdu+Wq
t/34h/ivGerR/mmUtUmQuIWgwCejc3uZH5CY8Ouq3cxERk0cwoz1E0f8gXD4TrSIvfI0qAYKxUTc
f87GH2zWPOJz/vazhMYcPjMnKmNeg6ddCHUWdrppv5RKMFotMlibpC07sMtV/OVmjVg++WQivit+
m9fsfT+ZmYwsTRmhMN2UutWtROzJJ692SRhPeWWu6dF+M7QWOFIf+UR7/W7ognUEmbC7xtnWNWkI
2RrKwLigMN8rGQvw4RAnMHeBOtM3tJyGEoe+h1FpRZQ5kTova4kgQA2TIksKiZKkfvtNEaZx0M/o
fwF7C0jvpFSLawxQCMu2P/XqcdMDtZEXx723UrNBGOR+2P5DI/1YCmPZWwB5JkVqha80KaeEfk2Z
xdGRIhyCd1FcrJ1qS5uXCHxeF4+aaoLwJvAUe1+HTzOClQpqyG9sEaOjY9XSpPsqmRNzbATCGA6Q
Bxj7aRTVypfgZDWNTmfgR+DaNYHTb6GiH0b/QUAeb8+dvna3UGR4OLCheBKJ0NyAFEfzvZtoWvk9
HmDi1SFcH7delKxJohXSV7Z2Gx371b4OIdOZEJuaoUDd8uKMxDiT67xz0YnVRZ+skjZMz1NIT72R
KQ35DKmzvMayGmQnc32jADoTgEcq580lunvWgxNCiD3kibw2+Dxqlx91Hrrw/XUbrGso8RBiqVxy
0eokn9Qp45bcs1yffJ+xER5WRma+ux4wjbSOQhhugMsqgPaeU7SDfQt8FZx+v8gvyZlwm0CWHVn/
U3ElIZMjP3V4I6hNNuK6JTNG2m+oSAkKhy7JrBH+oxFrEB5JJS3Mk5ov7ljQfuE5M3ed0j9vKgZb
3kgh88lnakjVbRmQjw0bd1Vd+7GoGSbyAma245IlhhVGXgQdwp5c8tCWME2v43DfZp1+8PIs3Ip/
uo9dSM6iOasPTkE0Q3NH0l4hCQR31ghzV+t7BDCF6pWbLvY8EyEw1Q7c6xrWqXyx8xh2sJezxltn
1Pq1M+0IQu0QJzbxcpxYR24EbAHJEmIIN7JJcF16Y9UasdxbzTxq3dos0Ggt3KRpODnUlnZ5vTtW
z7yHEPnKI7JDkou2HA8GQkhgFqxNustJQs8qC/dMTTvxmh82cL8UXhc3qvl0vdu9tB0d0Mu9SPhK
3zh+n7cXbk9Yu+CCY+NdGCqnqhT8dqXC/3YUHvQZtxiVsGqmT01jJD/3vXRGsg3YkihrbQ6muK6g
ygQd6p84/bW5Hi/jfIQqH8YvGWDonZNvndS2zLHq69gpnGW/22iWeIsM00gx7FM4fn8IeVOLt3Eq
mN5kvcIdFypXhRta/Is0F9CgOFCP8ll/Mb99vIdHj/S7nG9jgKDF9nxHXWw920NOjI9iDdYLPIld
Q2cwMJLufTg4Ljoxs15hXASHUsaI/g7NV0mxlkJMhBahYUVKz8jrEjFbNhxKLGl9hX990O7CWjCD
/e1vod+eOt8JaXdBrAnTynxZ3tgOnHyu4Qyqk6826lsHGiaogDtpNm5ZIvC2W9hNHrEDa2eB+aPU
SIFYq3L1TJOzNT1dPtmVjJpfxV1U4Ngn5AQCmD3BHY2fha7YPoAXuZsjYX5eOK/9AiKLPeZ2iXkq
16NALmEra557k0GqldUYxR53CDEv7+BYzZgOWCWmbSoD4F0IIsScvvBXwKwMsVV3j+hKHjKIbyTr
fa1vA9WDTNPlP2zdSX0sXleXj/4dpBm6deF+55g8ZJT/gGN7xVQNTEaoWnesJ7gvVLWT/UkWh6B0
MfAATx+jxajIoraTSB5TYzYo9y7lPOtzjMtqqn8+mnhR7typiYh9uuKqaPeq5OJa8i40b+KG5+A2
EGSTr0TCc7Ga+2L7XvYtGgymTEXpynOyliyT5zTUibh/MT7lY39ijFgeVvkdU9qe0SyqA0qPyxNJ
752iJ3FJ8k2bTYPrUmO/NpfgY3uRZhVG3kVSjEJl92W7xw9cuO6H3A0JveTHLoxDz2KwKRGlvmIj
I40CdRYVqcNeR34lqGvmF4dMZaACHOjvaU4HgS3UxCBR7DkDuncpZHPpcLBJNfeoYBpsHUFhP2LQ
j2gHwtTpsBFPoqCkFy+o++GChAoPNRvzRTqKqlrkfK8s5KTx5XbXKw3mF0SyAT+P1Ll9ZTXMyt3L
/plbapg2EVXg+SRXy+bAvG/tLmMUcr0tnpkIwhNKIahJumKi4vW9RgxERTPbI/BVMJnKpgfUgrqZ
CzDZDOFo3X3m+YP+rOskSyzLluE9ivWknrL3b8Zyx8p0tjEyhz//xboZ4bQ/+J/R8TgC+8z461cq
TwveSzq6vcmKPtyShjKxcLwN1vTgsZFs7+Cw2aKb4hOIe/Txi3oh5hc9ahjYiJ2DXboM392ATnEk
i90O02EpovFSWW6TJGH+K0S98GXJ6a05vF/w6krOn78EqYtcIefP6CvJ7C9K5hTpPElrO+H7PW8v
y0nhwYcSrXFPoG1KtsJEqzRoJn7nYf/RGaciHd9Y6kv3Ib2CZFb0JL9oZqaWJCGzHPEUoE/0Q7dk
HSi/5+DlawacIPMuvZ7JnvfbrARqJCZiz7Z5IHtkVxp9qdZKG0X6xxgPn/cmQEbu9AXMvrqPfSVq
Tz+pLds8gjVveXecVATl87fZBBBbl98KgZ/0o9OOnAQwkHd95ZnN70cmyYC5IxO/m/p36WW2KWJd
+iXOePrmIyM6aGR8t87I4D1AxfhvKKxmA0LaRjLrri3O+ZiqYJmhTvLpyCJa+EjGfYBEeyW4fHYU
Tp6udkg0PNIg4j1v4O6MXijyK/BErSWgkub+ReldTQ5RthHrT/n0LRx8nIi3ewjfZBhdq8rbvRsG
DxpR7CxuTOigPP/cLHSvGUDPaDAjBq+oNsv9NPeLJWCpgQ3aFuJH4Se4mISqCwi0IrnhOOO7ywP1
xDkk0p9mf0kSksLOwRByi+nJHvshzk38pQKkznLNhQnYLvTY4QMDA0DTaK0jMEjXxDx+Dh8lYMiP
MPKE+VXakt80xl4cpIBPDfEOhyrX0TZ/wk7vpkQWMx2+YV42B3TQsIEjSW+PFVPGMPankaGmT04B
Lp/POvOilG1nZbAm2bsUiyp+AnKBux64JCQIxQokA1BwvEIh4owFcMUfSYi7JbEX0d9Rqv7wjEcK
KSOgJXipBeFhLC1UKuSHlBzcx5I0eR4Ow9VeDvO2eWRnDIaRGWYxh1hQnhpgoSI/cFwho2zsQGQF
4zEbzrtzVsMNsEsh9HGRpMie3nM4IVl2zkcuveiS3gQRsbMMyP5dHWpoNg2Jw0NUSktmTLNmVJNe
342U887SiyVVtih891RgVb3iAsRcauXyttkum4zYEIOyYWuGldAhYEWxINYGKUli7k34NwbwZ70E
p8+MngPAXLvHfpsbkU5PeL13gTZuyx1YqQbMYMManhys/ZfzmbSg7rhWRoTSp66O87sbIRjKVy/W
LDn3RjNsJ0XJFso7OGKilpw5hvFEMu5rp51OLrnwqAOZSsfWMjwO96tsZdvxkR9EErC71g52Rh/U
ZtGVHqXgwwywECzxH2iSk6H7lGTKQxx+XcvJlKr4WYvTAfcoK2JLP/U6usOGxnG4G8TB57Mjizj2
mCy2fhBIpTG6YDpHbvxcNcSzJj3uft5AfRalc6/NBXnVuXFXMmNX5Id3qPENrw5/FdGxvfMZc8SU
06B4vRlRRSum0sDliHGYej0rYZIOzM5sSoo4jOSEqUS6AbxtdAZ1h+gTvlJsjtGtubTbotueZfHp
3yWcQiCH5BPSShGoHSNLSiKt2GmGUY/gOSTCcJoIs0yBCiTcrESTzKsxOkeF1fNOfV17xjjtANR6
bOue4eZyj8nECYzuTpDrZQrqe8F8DBaAF3QUIobX9En/jLcX0B8cH1HLnLczf+3OUKZ7UqiHNdhP
yqJx8EPwkmvXvpDAVgz313/c9Exh7eiHlWMQtD5ycHk63wMKlJiEbqw5FUz9S1aOAbOwc/EfGR3/
uj44xfkAlX2kvVd+7+XjaT4h1P+oM+t07j2bDXncMA/VJ3RdxdvcqroiYnG48IZ4M4fIVedIjcdV
NK0rC6DP1MEYETPhbqcD7g5VHTqGQTvQYsRJ9mX7Pdvv2DUv1G3Hf27aRjhp1GMQMfLYeWraal+6
IIHSp4aJePcwPKA/YffFot7Tt15J5jRtIwU3OaIodWetWlR09NOE6O8rY5HyGj6zBVjQHtdHCUZB
zhzxGTmFSJGcMmA4bpOhQzTdpnJVmUrOpNUzH87iGDf9HcPSNOc/f7g8bPhCfqRvOzJniszEEVsQ
3RqCT2Ni9OU/nwURArM6xr2O1JbpIN1Ew/A0I/wD7jfmyqcj7Wa2oytCFrPp0/tPdhNXJ9L9uJ0e
ohs344tOG9h7drEawtcLYXCpn8W+DvboIvKUrzcaxFO3vgWMTlSOHe3XN1CH4+8Om1uo5XBPgt/s
YP1bPya7DV+qTaWD5KDuVXLEDyKCJUdXl0IMHXFF7vzKrx1GqZ/viH5InZzIti0YV5amPuorHjjO
+0RsplIkT58/YnWQpc3kCSBJpcs142IdBGgmzRNYvYeIMQEtTgtnztKDT8hHsytWpl6px89GRJNp
Z7xehvFPkToSQ2w8lwCcLQ2xncnxNEAwvsN8gFbseeJ4Eux6bCuIYHMgFoOJbJk05/SAMfK0Zulz
U4HSDeRElU0i93i52w3pO1cZMjBuH8tQJphA40vuj3JIKaXtDt3WrOL+MFwmf+cd4emYoU3B/ONN
/ALRvYWl5QpSj3318DV+559cITdNBkqNFkUZ8A/n4vChIviiSi74rf5/4Edqo1ulDZS09DtkpisR
+vswzr4M0G8P0M8yeNCwT02Gl+gWPMxdKK+SV3aE3Jb19d+hRy/wImcgj0Bxmx/by+jma/I26C2m
Nkt5lEFY2wi7cvh7+4JLrX1g2TfnoHJhMFGLDXDJhhxXP9iFgg1MH063qlK7OyobFk1OGj01IdDW
IhqLs5A213+CRro3mm+7sLGIhk6xo8l/K/DZ2LhuQeQ+7aXhw9psdRL9zXoy61NVhVajxCYmvRKF
TqXoZuULI/JvxWuuHU0MJaNqW/mwZtCz1uVCVY6jSzN8mFkDvmpBtL2qyGu/862YXLS2nFb06AYH
ZY3nPbWIFP4eXcPK+KvZ62hCLvHLH8KB+9IneWXZqGrqZ0fAkP86TvoE0fy3P0dEChnKWhenUxf9
EDsaANw+s8zIODMK/N/Qbq/qUIv7VD8aK0+V+uID9Awg0nS7puY1Ws9YeaIUz0ycH59eyyhmxlTg
y2Jq1lLActKi0hdbQsMkV4BLizwnybq+EqSXJL+xU6taZwXftA8DeNn0ZmIyxbkk6ae4eafHQaO7
ZJdjiv59r+S+fmmUuOPok4wGsWZgONLBl5gKW3eucjj0KdzjYaPcALmBc8y1oPQb5xyObpeuox3k
8RRQiGZZBwbJPMBUjVj1cEWjEvUPXFB3vQQFNRCMHURF4i7BkTp2dbYplA+CHqN0t0LM8vEvVMfq
wSscXTliAYP4yitkIF3aycNGbJKP3L8dITHtO1Pm+8aLa2Wx8gjsn1CeoQVlIxJXR6hjKzUoHxFC
2GmMUmJyF4N8pFiH7MHAni+e3ZnBLTN9HBN84WVAnCQTrjzOe6kfy+ymEIGzGUzB6wK/zJuDLATI
zObwz0Jhyveae6W0iZgwnl+ynAt728ka3AIsKti9ZKdmt7OzuV1OJbAkR2PD7snZnxP4DhO2ADaC
hKAiiN7RUuvdbQeoHBR2CfFy0W9nNQXyzsaaDBuC/HZhnsUhCKrRXd9pUdXmSuHZ1RRv/aRKN4ge
T4wAWl6GPGt368ufdcEeIVre25EFFtm7CgRoC+A+kTO2/xLI06MmOY0cp3NLPn4dJm1LwNyUny5d
EwiSw+NYc/0Pi4msc5An0qOyJVaWuYnUT4buALWXsBcQ5DTfbk9TYeIUrGLfCa4nAIW+JYs4G9vH
+bFsvR88lAMkFvn6ucLZI/r4D0rEiem1lwgnlNbiF6AfozfrKHYE1HG4rcajU9ttjVE7Uo4l1wWb
aLvUN0OVM+c2Qof6Zdtk5OGzzBd2KaLIFQdTlZ6NKd4SfEQWlTQKWOz/1T0yrlfwTuXKTneAwkhT
rqq0gXVA+ZeDe+/sD4R+3j4gaWzIkjb4HwN2YvBmwR9bTEMGek556sMG+MH84MQ3HH+0KvzO2ZGM
lIp/IHeKbqpUpxuqN/d94vSQtGZGdtY883xUaot1bm4UyEqJjoltqCZMIi8oAY6ONuikmruUTYo1
0A7GKsu2FNhEpo4/QX2zIOQI+WCYtP03GsPykTmQqFLITG8k+FmQN0iyribQyL1dmvSKAscM/8TU
cGT8Ecxrh/Dp0Yf2qKGJL7Z0A/DsZb9mg2pjs+hFLl8Tc/MvydgEL04+0SKFVmOPYJUqvtYODHP3
YAwLMJ5PsI6fJt/LWsTv4Un4xiCIzR/IUZmz8pqc0EChehoSW8Gt2PrKCY3QBazrSqh/cO/e2y3A
tKgmKXymbfpYms2N2GGgzpFlqS+PT+wnXazyUoQwTkGIN891eTWak2xXKLSZJx9i3iP2JQ9TirFt
+IZS8y4UwGRpSu6xe2p6RetlhVpT5lk2X2v3sl3ZKrbdqvgV2IlnDPOFz3AxLO8CdmH9g/oVUQgj
w5HZydWXqL1vpzUcORxKMPo7Z+cZnIQfosWsYaSIP0h+TZD0g2s4eSissvDMWtAL6qhckcxvKTYY
ud6EuFwupeneFvoKQkUyEGIyQ2gpzHi55eisASAnoJAzu2g9DtnEDJnkiNldABD0FmYXB59oZjZk
txAcvXjZ7iSkT5hcdfkcWTJI6GYx/ysD2GR4d6rl7VLLRTJYcnVbuNbFWbpEcdMQyvEiS0hSsCRJ
QhS6zO8iL218wWW0EbjcZfXHpoPoZCGyUVRCv4jU+I5MCMTKuP6H3TclSp95z//pQql+o2Wb9vYH
reNtEski1bAEdYrfvI0aPcN5xJUqZM63+bHCF+hb144MpJMepNyXU0S+dUYooHRhNCWjFih9Xy/p
cWidt9JK/GBz5ePtIW+cnZlKYY+sUPzaKE+/Cp5uYTxVJM4bqNOzNeCKrNar5ikpv7zVKXA4UgK0
7AzZetq1Yill21nWud4XcuFBY4fTIPrmdUHFcpGrszBKujEwyiPcOlwsd2sS0jg91PEOfzNu+mEa
JHwSjHIKKdW4e8glXFnt6ppMrp7yKDmDfkRaB6k8eQrdqJXOPsXosoBrLdwAugb39Eh7GV4OVUFj
U/Lw31DKCerc7VMsBnlIrBpzx8BOTXVel4WLziiy18+bOrUsBkZc5aFLMlYVlLYAXCrlw/isX64N
tq88/2rR728kpLjR02S5LGrxM6ApVsoQrA2JgD+/ecIR2FyNojroJyyUJFA8p1uaNcr8veULbi4i
7drRthtRPwuU2RscgNAqw0pP6A7VZJDLyEVf+pX50WyQtYBnKNkMJ4FZiE86Dyl+EW7z1VDM//cA
hzws8VWCiIj3elIE0uZzyso+Dficip8aNLtN30Y0MrxXkd3DHqbPRUCxMWnSt0/cyV2lbTHlgXNt
PAWY64YqKo5CGBpS25VkwAoHxuYNqThJ63xITssO69gwT77nbPipek92KJIBLjatn5WJRue3d1EE
RK2Cd2mgse4rnRm5xdHpapOBn8M3TWS4b9Rzji2XkxtOlRwLEAIoMwYBZFJUStPQh1H9dy8yRRsn
Q2/78xi80QHNzEcW8+BLcV3df1G01/3XZAMFLtPnmm9YXgTQ0AbQT2yOiAucfm1YCgO4if5WGis6
k0t+4XC0KkoieZJRyCw5W+oQ0m5GMzstrJJ99rQPVb7mvXnvl/uRGL1VhQ5r1+FdI79YveowlGGU
Y5kl+McE/gcmTuMl4UvrKDQmwRRozqd33bcHetDe9lbP/UTim6SbpIlMQhoKDP3YRWDUPkH9riFl
B1hUJGqVEn6LdUi/D19ZqZoh4blVZzH80KwGpsNUsfJHgz9fIH5jBsJ8wKhrZI5cPm1mjdT6T7nZ
zhQ5XZ+MxjqmUhhZpNlhOXDuL1FlXP42dJXtxm+CIdv5zi3KUgrpdt46uACLV+SqBm+ySFQrBmA4
oMEsXTln/TJ9xOWS4mGG/MdLiDs+nLYaXA1t792/qptaWrgSULMVnHFgae+gyhHzwXY1aIyRr9OJ
CwNsBN1W4Xs2ttAQCt00eNf8iKlsrP0luvbcv2FSm/Nnuot1AuFp4p4hprh3lO0K4XI/gdAJAsJh
O/UGCxrBSj30rirc3oQMJ2TFPh32IfDVtHVtPiFwLYvujVrxqC5iCe+2rTS51JutIwh/RBg75rqv
JZT9jf7gqZAFt++HtFp/1Mk3ZPlJ0vhj71kbatEo9DEQgGOgpUGBpayDIZUoW9v8v8qgkrs8qGQX
v7HpRjGYzalm7hEFOoqGHz0/KzzEEshfBwUPvkP0nwDt1nsD7QeNJSQDHw+T95GTVZJlZ+6nFtP/
jHZ6HcEv6wU75xb2QqA7MRgG4Zm79l0qpjsdtRydOwC2iItRlwd9NNk7lfAJbtNF9dxD57z3nVn1
nG7g2XfyncL1OBaC10LqxxeO0ui5zJ9Y2MoqwRY20SdifJqAPkLAHqjzhvH+KCEkzCjbw6fsr2pf
edwdDH/4GIpeuCPGj/cZZX6o+iG6rQ3Qv24HfIL79ed52YIvq44nNNweS6KIriJ1x6vCaPawCZXW
BUCgIGPLaZsXwvBUOszb57mnjv2ACyX2Fjw80BohK1K/748yeYa/aCusrCONCPELSBIuPyLa5/e9
lIPVgSTz1WpsShzeQrSLo/aq/jsYfgmwwTgM1z6w/2wxcSvsgf4CTJO27kowZvWXbEetd3822z+G
5uKSUOzFKuko3gZGMmEP3o/LY+TrngXugAvRDZHsXBYhvsV+Z58JZsTujQdRSHfCSXfNDHQihzrr
RVzBooxtD1A6UtMkzAK9OflZpQT2cTS/98X4JMUhMrE3VA9cPatEkqvjmT7Dxwzcw5eTUCGoOYOV
Gugce/glLv5YepEMIvxy1SLC3ilP1bbcOYVOlZKWicTzrb/YG2zEcGdLsJJtfwCsWlCqgJVrVsk5
gJX/Jzs/7hWpSyYbWLQYkthjgIJkiWucpLfJ+a2dwqw4iG2iLNoGUk0LsySAjhqSAbmNgdfKGa/8
PVPSVnlxgpH1dxxkVM65JEKbwprz9jAZ1dgjINFFfiRxZm+4Am2iHR7Qlphh7BSOAP+3UDQUsPz+
0Hl07gEnDM3yEJjbjtBtzGAHhASOJ6hKrSkq4C0+DkxZveLOA118b9Uj1BF51G+V5pLz/p1oMAOQ
YdirpzuRGQnq1rKidCbzbRlUczZomazIzT/9LZNpnVqxG7PpiO/e2wfok/cw/2CTZ9BKwedzwD1O
3ernjq/ZUoO1GBq4der0nUiYc9hHW7bSmnTbhdcYbohU6SJGFMDbqRCsUqtPpXK/qfI/2QEMUtlT
m4p27sZy4g7O9oTWp7w2LhdUG1AG8/uROHILUbcmr3fm3ez5inI6kCM9HSk1AD2TF+j46D/21ToE
zHO9KvywEWAeyjdqVFUyous/aSfVd0pw+FmW9WKkyJCBWY7O25T3rKn785yZCIRzeFD4pAx8qM2o
yH2r2c6vCVT/GIsgF+cHxHf4JLkY+GT7ucWRd8I4bcMnE7ZW3xvPxKUIpajcUr42c52MUJ6Y4XKH
f4+bHmyE6QSBQESJXwmkRkxjcjrR8k3I5dDSTHswy0UJ79mtw8W6imJ5221dmdNmQg1eqtUcciB0
MlKpk2Pp62eFin6uy7O7Gi0uRuxT6BUTz7pZjuhKaBW9h59orQIG9EHCHg9JwCaOIZBELpA9zMzj
Geyq/K1t2lR1Od/add/oW4pX8xUTo27+NRNkz6W6e1iO6TgMHftmG4FMQGUSeTX8c82cRlXuu5uE
CHKX+sIJyPGYYt5h93sYVWNw7HU9xQJjhmIR8u9OWWw5tf0ObO/NnutsTYifbtO1fhmG4tup7Kbb
6fN47lkTPvQU+U5sW3LXpYFi/PJ1a2rw4/H/hqdrg6ZhE1pYmX1hyiNRzBrWdPQ3qoEr6okpE7nI
J1DWBdAAyeFgVUEW7CoQ6Px6S6TtdyJlSnzLiGQ5KSK88JU1VC+3ktETtcnOB6WiiIKpz53sJQyq
eQEJ1OJbP3cYBPaTEggpKX3Fe0e3MGR69f69jzaSTYwt2VWLin9dQBwHhK8is/3qrz+shKdbOPuQ
btiZkGk4lnIKeYwAs3J/TM+jAYRHLxkCzFjh+lzmG8EGhoqg5VNC/TQWFgH63uAYa3kvhqbBfaGz
EThG3JAMfG1b0HZh+Rv43/jtdOblPkbhgVykY8HxAs/Xnp1WsmDLMP8s/Wd5H5nyKr6MSDjyJffP
bSh+L07yXahmqSbG12bmIR98rteJLhOjaJFxw5iihaCTEiNNFm5w6G7V8CZIvwI50TkCgkvLxleY
AMHNXRFUqyrG7jnUcAa/DVOqDsGfnGaZD3S0mbdidpTq2TB9TioZayKwq5RCRmG1oM+2DwxkuafX
gNM3cbTWDmM7HBzIlB7glFIcdzyNWvNjgu5yDH2vd8WYAGmqS7LqxijTXOwSEahs2Aq+6g4XvXug
u5tzzrl34Phs0Un/IlQ4MKt5woiHa+2Eo5nYMFBHuTBHiaTCSqMKmUnoS++KFtkd+EmmqTyXpW3Z
pC1m3NQ59rJb+89U9mK05q4U+VmjLft4yvcrzRKxcglGw8lFkFdBnirbsPG0Oig962S4C3uE8dN6
Hw/na0+i1OJTOJBPbPcGQ+I+ZLpnklaaRoX80nYdHNSju8vRJAT9+hBl/Djhursi38bofLnoWvFy
XqiwwI+R9DzOJKuR8japPpaSr6yVL3eMRN4lIwS0ze25OSfQc+Vpf/4sd/EyNJkGeUJ4bgydp3V/
QoFSeP0OrsEy5NW+dBmmBcnMsfqNO5noVetov9v0YjMfWV1Z1DdDF2oeorOwzd3siavv9xncJ29Q
GW4cZtsOzU1oPsQe9n+dCHjxyACD18TK+fGvPmsnKGSH78Tg7ubQg0VRgsbYVUzt0U1VlC8sP0sX
gieRB89rvzY5WbaOCXtl7L1jNagiX6irhXMLOLeI9QO9z+8CfMbJ349MzZTbI4bZB8/ZCc3Oa+gr
1aM3ZB1z3s4WiljaNpiLUl3d8pKXdkKV19CUlZrTGF43/K7LCA6lr4e84KjWJiyIz+DipmpWy4SM
iqimuC61rpXe5kdmFivttUMQDfMV3bSqLRklc7ud0JuGdw5yGd/L0sHRXElj4081llR7dFNdq/95
naGh7aWwSAeHfvKM2Wd6tf53N8jLr2e0hzW51Kh4OxE+Y12IH9nY5vZf+fm8OZBp8sYnY7PIdT0g
MRr02jW2zzLjgDZsS7OzYcCJ0fBfw1wE/GcOzBPOL1yUQvLOrvXq3XIDMfkx1tpUuoSvstQqp+YC
FMlTXIN9zXhOw6bImubOl0FvV4ER3fUhhFub0e8vHg24mAyByy6X53iuOtrzC9ZlJxZTDN+fKhXN
IfTIlJcJZc5ZKPhS83kIu1Sv/joG2Di/1l/a/mpagGKTW2x0iDCXzwyzAOtJgKJYu3qvLf+TABAO
SWBWDGEEHNSuepRCD2v+/fcpb8OXgCdWvwJBCMW58wKHB3+SyXrBd8MKSQbQNuMoWviyVO1vDhd6
AjwGdtGc4GMkOU1L9wPqghzfJ+pY4GKrshD2p9JbcWxVTdRS6ShAflBIqFDow8Ly2+7IaQBeWYmY
qeb5nEVADGhxFde23+9H09qrUh0hIFdMhNU1JOdasmO8rsiVZ/0PXnU+6AgFL5dJksQKjwhfTyyt
vvkT91geh5n96e8F4HPpUwNFJqABnQ/MScXIpBeR/k9Sk/f0lDzQJj5HcV9IInCG906q/y0kQN6n
mBRSokEd983q2J68IlKyrkMo/vbR3qRBpg/pFVo7V0NuBHmW/OqciWRcwvSerONLDKEzEHdl/mE0
Mnd71i1APSPLPiB7qo0n1CH7AcqJPt5qPRMyuuiDacE37UvQ9dSbfICXQyyok+JScmkysjBG/C/p
10ZvNZSoIFLVWT13t9gj0QG+jfeTdcNuCQdfUDPyaBdJ78htsZqeSEQLzc4tkat3XJOpM6LCioiA
macPFzoI4GuJpVLyPWe3EcH9JZ0J6hEGTQdHF/7s98ttN42Uj6127oPEddz0uVJeb4CgWTMibPa2
2fbbbC9UgAM1GK3NWQT+dY4v+uoeo0NnxSrnQnSATM83PHjlkosGVT9axwvr7wdRzwIzp0wK+206
gVtYEkaHchioFYgS/61JKDyHi+EMDBJeqOt9h9NQpfi6l9GR+DZmyY95LhbQ4rtSZe0YZPrt2bam
MxMk/e2Vm2DX0wkPDMFy0Hd9IcbJkpubRrw3EdgdUO6YhJPpbRE/rXMdSP3OYlbA6wMN01ps8f0C
62eB9NIL/7iet0cSzPnsOsJ6dXZU5cCf1DEdqUJRpTOEo9y6BTyH2iZrw9uYy3mgvItQZz8Gw12+
icSq0y8zo8COHGBMoY9LyPYA0McGF8s2y1ESgtnzfZk2suyJQXSXxF5nDsI0uM663jwMxYzwrBhh
5upysnv5N/6ZBbEQrcqNEPtxCTszjNCcT7FgfFuuQX7B7ZglRQQRrzYfwNgsDv8DevJuCDnGP4xq
XPB1h4DbU1KquWDGO4mgNuZlj5rYuZH/BiY6LYHYRdp8csK1eKJ2QuYFMv9jfhXAeSCkOHEHzj9X
bLZe9/mOu3kbRGLN3RKoz3djXgIBeigSi45PORazBFCqFamPkcDmFGvs/YSLN48tHBugGDyYDwit
kVbtev+fgUqJwJaBfNUpTR04I0ohRdpRck70RAU1IS81hypkzOuQdpcOVQeUOBaSfBNFbk+vEYUi
AL+RcOGdSl+W28xnLVTrA9jyTU4uBZsMrUHM1XOM44bSWJiZCBR0rCV/FSS7wQMT9cJRau+TAGS1
dMNsT5huFjZXfSNGepDw64qJIqxeRFJgGtY1B2Bw7bDI5loF8bAHQxIGiX0S6AP4LXeojlWFKrvW
vymUFVqJ/1OXzyUh+wOBt+F+Btd+RqEFOGwVetsPWdMkeXXSx7NOdPRDPd2SYbouFwfBf2SQDWbT
f+xzov05I0R63SIWKcOW6AG4btpm2ZY9UIhOF5xbBxoiCPkhTU462CHiK0Dl9evctd4dqvjsS5iH
0ZQGpQm9pCpu5LzrVuNo387uVEkrMviyVU2zlKUPTL4p+0ntVZ+H24sAcVHJUgJSAdF97bAvRZbg
3ixTU4MFyd6I/slxj0ZnhOGYuXtxIFfGd3qd5kSMOoIAyH229Rc7nlRRSmyqj0mT5Huu098Zxcgh
8GjwEHEsuI80wZDLjdY3aBVYOOKw+xqjMH3PpE/a8GI8K2v7NHk4yHtavFRnnL30sjn4SHt27RIT
6AKS/qv1P6oNznIx+lYm0tQgMBUtwd325Bo7v2xPbh1I6N+XKtCjxYfqVi7xm8xDwWK6VhvhgeOT
IU4TodHr86PmE0YwKHndEpi+8Jmhns/NS5mdRLp5voasjg3TmFWoKzfVIkQlKi5BxJ7FvFJfrFGc
Thb0nTGQTYPymGGE1G42u8vUhGxhIUNxERkwKAyC7kpRIte84Hdtuxbd7qlsLeqZfBf7LWqZI7eh
F6pHeQGxfwEEFkiHB3DSl8Bmdn/bN66mholmAX+Pus2K/xvYzWMaIbLIYlWuykmvO9xUHLbD4tuI
2wd0FSNvAYgSy1uXbmIUZQ5VcKCppWarOkeC3Z9V/k2+9bNAPjQ4AKIUN7OvH4dZe2LNMXgIthoQ
S2LUvrrOZuQ7bqVAaTzXpj3E2FkYErBHN9G/JWz5Kr+u3BWZOKU0pkMi3GFRQyXYBkPFK5ku+eQg
a2vr4HrqoNVa9UuWlEhuYXMG8VYNCq6xi3Q7zwqUdavAsGfqLzcNCJs2u/GeaogbHCKumphMzHKY
7Lgi2L5JjtoczG//9yfjxDa0qdGmk2MvHgZJS3HYv5CHJqAt59Uc+fKoI7hy8eOOgxiNRl0G/16U
wmA/bRS6P3ayK9OFR0zFJKcnQAeSDiJY8VHptt1AlDTVmnDKkZS0D6Usq84Zu47uarsCnbOn+8TV
kCKCi8GrfJBPNl/scnORGEqQR6hjVZNNB3bI7fN3pHZgsVY7HiaKPNWcgABe0QvdmhIeeaGUUNPh
e0qFusIV64rjlF3oNaqCo5+H7KkxGhCdRv4ozoDdLXtiVoEwEOCdN+oSQ5loIj+Z37/cZ9AxVgJb
cjlXMzf1UPD+8SfZSg9NY+0DEVxJwtd23Jtuu38bF6m+2flFVPlUG0jMEwqZGhbkOgGxEInob1eV
qFukDzMDh0T56SOzYjIXCRMtNlUhF4TNRDvJh4fYz1SjAN37e5N+kubDfloVr1GpLGiuuvfvJFRL
/tivjbZgmeyBvWaiEgzk7eTwxHpqsEB4BAl3UaU3NtSLunQGHfyTvqYURFX3jEjcFVWh5no4K1P0
9QV90JVoSLtQknOkRxRJx+UneweilbysreAItw8IQUazXm/y+/QorYh0kCaOxFcM+CiaN2a7MpDr
AAHLc+D4qPJPcslNC80oLyMp5hAMBXeObpNg/GVxHWdNUYwwyykYfUuG9SQMzY3jsQEV33Pv6Ryw
fGXhwy33/Cpr+0IEOqKQmPCykp6WD90YaB1nhaWbm15Ay/itK7QrEOxgCNS1E8cEwAWSq4SBVIb4
ALvt1LK4Ol62dzC7CJRc7zYM88FkkCem1eRmLN4eyROTEh21oQlR17Q+iPRV0+4s33FgTfM/1nQr
IFQnbNmzvgNkP48u1G/xFY+IvpK/YuhVQBijuQTDIWLlr0OJUFxTYPuBRY8Hv7jqwlwwCslUKfsF
SQdrey+rFLqPErnZJnLv8uPpdas77rW93r9T4SggP3BAWhOIN3cboBCWv8TvUqqx90lbLYLl0LpQ
5usCfF0ZlNkzVISCd3HfZ+bmQIsQ/ILttJ5OugPj6c49KFORDT4j4nJwoGdmTXXafqSaZ07j6HKc
OvCCH50qi7Z4tuRwRw5S4kzpm2jXqEPqVWtRoFTc0F/i2OSxSKrI6eAODO8/ujI95XeKxbNDA54t
WNgcAcyp2fVFCjPGOtA9/a5Jt+bTEayZxOu5f7ex0+l23fFcXXgySpYoFu2iaPIPpIvo9dYOiY+f
qjjPsdeEPMNKO95Waq7VB/IgahEW2XCJz9ZN0s1EZjj8iKfck8Te4PbktnUUo/w+DUZG62f24ddx
QWxvI2Lt6q0aM2zQTmCc/FkxlLwjwRS7sg/2Ow+vznEeHOTwLO15gY2KYVG30AXSCPOtnUWZAze9
d3QzJYJZsTAZ/OwvZEU0jahHSgS4vRY8lf1MCtDxniZnLsyry97oOJSzoY7Md947C4oRT+Zm8A7z
S1zdCDSN+4V+nZ1yGQFBVtamTjQoMWt2uW5ibtl6DjeTw34BSayP+SrWYHYUNoKOAc132yh1Wqi3
EfM22Q/lESun8Zx6NsPCQKmMgC/T8X9rVZ7v3Rv6MRs/sYmvj0uLbZ7hg4XEl4p5jDjlYXgf9WHt
W+gxfdztpu9jYLL9aLC2M+h3QO3v6q+2H9qG61/eJMKXIhMGPiJNXpFiQzoD/gD9XSaEA5oanHHk
3sJ6r2Ya8G1ESRDbZg2srro7wdVKZ8lq7GoRO8RXnAQABOEpMw/HW6xmTxNPXO2dd/FLwIgsZWdy
KSINDpP4sG6tou8GaOoRKqGU3rLc8KNcemcWRTxWdfGSU4+eY3alp/1cy8yL3zZsEsnf9tWI7myo
mCdkpAw04B2JS13OS/Prs71b4KOIod5bz+e1qZ4q/2+h47ZHi3FIpzXLmbX7+x6NELIIFgjiVCu0
cuuUV9P6nwIrRgjl74JATHqW3lj6Bp4PWKi67Iaj/VBI36OqlywKECdYB18zErqC3yo+QX/W0ZSS
fP1tysZ//z1h/eu2+AEbPLxAmR9Z73tnFZuQyzULttuXlHzIi6/VzPnbHjAs+Yis9zLHqVe55IpC
7tMl4uKlY6DL5QqARZgy58BbZNRQ0K7E2P6vRjRN5Se3T+UWPKzrmI8uDOObXHbCV7J/QEsxvNhp
xGtaqbxLxJjQ0EWlMeJprrNeb1AcxtBknuhnjyolUEVPoSVlII9DaMc2GbjueQlSE3F2GlarMHGT
RvYnAYYncsQKJMUnDyO2Ujc8QYzf2QDeA//cYWGoSHpzIZFMr8KUb4AuXR7sgCkilue7ejwUXsCm
oG9I86TxZMfOCMjKLya8TZxa5HXxqhT6hGQLVKTocAvSOcT/rpdpM7uQi9HtAQTfZeSlHxSprEgI
2zqern1poN+aVoyfcOFUIexqt85MPFM7jonuouVai908VEuZdbdLl7lRdXHTAPbAfemZC/Ks7g+G
geBIpM+u9sEfUQR2xY1k9b9aFx1HOrC+VlcHiRdmj03/97A1rZ5JwJKlMtNzgdZYZVE7Uiz2gJLy
hblYidH6WPEd1TuKw6V0BP6optGA+tcQhFvDdfei4P09nTpTQprGCaeYz8r8GS0Y76vZ7VBV8RDr
TPX41mFmG4Uh5Y+btaJkpkDLTKTKV0nnK5E/DTOSWx6hhqYsi9M9fLqgIWSVFbk33UTiwTMRG+H1
TQb4BPYVzmZdy04+k9SRiS61dsGeJcKdTUN393xqFnvDzd6uHGbBxkWym1V6bgc3C516oeGYc+59
3crcxPdM7Xa+2mdN1ypMTXxmXsCSldup/KqTFN08AqOkpKIG0o753BRqSoVFRtcdXCzvTWKSxDCH
IGts4vNKDBoYLgGZlXEowpA4MGpaWzyS3DyE5FIFBGiPMIwe+3vYzAO0QadmA4JmS0DF3HerysvD
BZxsVhaqpGRhmcEbr/ZcCRBE45E3wviWIRwpI6VczD9ngs7ia2wBfLBxKpnDBsrkeU3g8CNAwApz
Y7e/3YYaU3apvFqss735NJapK3UcQ2yjFtBTgvTffsLGM/8a31FyRgNuleZkyqIvIE8hryu5l+cD
81+znNlgcCmwr5EC0s/MzwPFEHoLCGiu9O2bTO9NJBm1brxVyuCvxLIE+StKHoW301W6MwTfUak/
S0oOa9RQGkYBZFOhe1zxbiISGi+l+cnEGB9yc5sUs99sVpPAh7mdqiFYgNtNKOj3+rZS6y4biClW
3u0XEvcPjXfGnXnaL+/bgIplIil3/UtKE+31bq4DIzMLWzNPiI6RjWkJ2Dkv3BLED/XIrlsK5pPZ
+9rzw847bfexOHjq7HtMywc7pxOXxiGIjxP+FYKBxfbAVXWOdC0IBHT905D7HzSYJsBGmRn9bQs0
KZyBrw+NAR0K+rJmDzOHsnAU7HgQuBdKiMBOo6IX54xooe9I+6qscHJZ7Ug4kuR/9+dhWKNLR2vw
VxIpCEUxn2Vj/zkjP5ks07U5bxWWy/oF34jndMA31kv/29iT/ivJ1GjSnvYuQIOS4tXXfYKtNUoa
HkEs8omroL+proXXThYfYhB+5Iwk3FYOjMVmALFIMKrpPW4eTCTq6UKXLhPVdxiLklE+P8gTbpYf
9WjbCH6MU7FnVRbDXSvL7MneKb+TukaHHNELOR8x2x+oQqr7exPNF8mW7F5jmrsKYHbDcnFuKdLu
YomhquiKcPlQX9pS/MRHiBkpBiEFYjaaQ1156WJQLBgh6fBpbJPzWmB0WIpkdtokSwfb/VnzmKXI
0rAcvgS/nRcXcOdHlFnvSP9qTaFni2gO2wgTSoT+A2crxUKWfndyXd3VXX426T4MKdyiiFSKHfw3
vp38OPvPlOoxKF8lcAULIExMcGYrsXakzHP2dansK+8G0KmS+kQaxA4mAUk876JpWWDsAxqbG6wn
InVhJLdZwRI+LqOqofKM44mKK2HK7au3YBvDPzMXf4Swix0zb29yfssSf+GpyRyh030/Q6DY/GS5
xomG0GHknUAoBUcRTzWLEvlmgwEKZek85r6rtE2wKjhLixMumXRPtG2txZUc8zVVpfpQLfYR/U9m
yV2ITQBR6HXA/byuymnCkXv3YVtA1EouB0R8HDAoJwXCKYHjqnTcC9u4Vv88WonGnDyn0mErl3Zo
isgA9nLZvHJ5V8d1Ndfg3l7Bf5eA0Xtni3KK8g2//smr6ElaBaLmyt0bX745i8lIlv/VpkgavdNY
HbOJurtvA5YInqK8rO860fvra0YtDYwf3ITp/Mjs9qcKxdGjBcp1TBiw3r+f3vqoblLLwyISAK9U
ICTBBskb751vTwqdHDOTUK+Pea4GUSAnT9HY18wwz1BXEjhCawhVf/dj0yAbO5aPjw+UWfLXjQ/u
r9dpBorhYR/LE7OypyTx6mMGsOfEnWNlaXhDNAvJdAWlPY75mTwVhUJLjxPwBuFsjYhIT0ikPp9u
lFep5DEYu5j7PD54ssIFAaL8ACWzLlmZrxzp24tWZU+s+yNAgW0zq4KxtaNh3w+5u8HxKNqxDWsN
4vTGTgwGrMjnKTYYkBFj+GRrlZq/3J2gIqihljyjesR9sRHSR5aXXv9SjXG71Hm7rJALHRlFl9YQ
DmQnzAvbe298dd5fFRH1es6N0B17SZ95M0vl+DVL+V3H0vOQTeA/Jfl3FXkA//lSpmYCZNdF6Ij7
gZVo30i1K/yg/fooRF2oH3Bw8+3jH3QygnIXuWaYAWKCeY+Jn0+v4fHOkCcx8em4vq0SO2C7e/Ei
DUORI94X8moJpDkgC2b/xcS2H48EEWdB8zsvxlo9qrl0BcyWlXcTvExE1pFgOUWDOSi7Y+LpYNoK
lhFl3cddkXiIHwYoDEyQ6hXaoVE//nophI1E6fk5qu8SGczBwpIc84KtpuGxWK8w12LrmMdN6eqR
s481WW1ryxwk0MIXEF4C9WOnyutyZgejnoxJY0nu9CQCMrYquER2WW5iTJXoHpbfQ4nNM2N2bk0O
INioxUSDMOXFL1ZNbhP168HhwMOHkgZ7FIFReGcP5Vd7WYwxZ4XUV4Q1vFu8x8M2HCivaOlo2Q+M
NYScEGZ7vCM6OAzujxpH6IneFLElysCbLxHTeelhhgl54VF0myyEFwKUdTgzWFXBJtkVvdHptvbE
SMg79tjyux42AkOl7Gc3W5yZVwwQmpRHQR6JL4YoQqdJJzfExXEtGlwD9kncctsR4HQ7EO4j6INR
ECrODiV+FVhfSzCzUQhRIHRaxmh0I9QF73B3Mq35qTPFJgXlIJ4olJDCcwjIGx6k7vXijKYJhPIX
7jRbRBdRp1lTP/EV/iB0H8FtEDoVaCmlscHTNVM64F0/fyIXo8DxWhPJeetAJwYUVnMiNdtl1yVT
HPy/ItMUtatIY3He2SnYP+zFKA9WSAo7gY29WOivkPm3AvoCsMRoYCJyGOQW7BJF/2xwNyIW+Pvu
BOU3Q1yJPujRY4oT4rAWzf8g3e89Gwd49p2WxEAhd4yKGTP301jc67Ns++Mk44mVAOIAqREPEouw
rB3MSTDhh9Eqlan4TdhEk39jaIlUjo51XVnZFYwLKV6ybkIb9nfu8YZuffWWpO0o8X7eKm6NJfvK
2Su+dKAEs+gLLZPCgtDJpHwASEupkz8jv+6Z42XoJZZQtnaVRyKKOqTrlsUXTcQGEUAjAfeKL05i
027I/p38JOYKsHznsy3TMkEObdj7dO0ttvtq4akM5bz8msoRqD5Q0KEg2Zj/roUrS8rWnDwX5okQ
LreaXgLT8k80Xvw3VCMqRcO5oIyiBOGsWyLW3LOZOpTFcImyVVwBHEVouLsD3zKpsraHKZ4pWOMW
UCwipC7oTw6DdDGKfbg2vTrGwM6dLp/mTym0vmj3AA35KBBA/nhUpeIZKr32qYy/4HcyXQNVLr9k
Wxc4fTt9PakWyM4W1X6vT2WgYehbBFF06J27rt+qliErm7wDgWja+prCgnEGaOWDtu/jpwJ4NZ3Y
t39eWJV5S6il5r9/xdCWI6cWBWX3jaGfR04TARtajBpNyK9WxebqQCrhviyfWmhynAiED7kyP3xP
hyjc1PWcu+659oV5JhPH5YkRE/pXhd7UChvIIJD3Rjs9f+7Z/GosF0frkeqF0/K57WOT5QXGUmK7
h7TOX+RNAcGoZXasC98UpJkp53ONLpK5+Kl7UAI8tzKZbskt9wi6dfhSDlNU3XqQwyv25/bH2Zs/
DAnir3sAV/2CeYEXGXaAhQSx6QEvG2CYzCSelOY3Vm1L5EUvIpOWG78UrfQ9zJhZEGZOhYQMj7I8
U2xHccYREENEIfzrhYwkD/NKkMaBxyYQqAjCYeChM8yhGHMwGwZ6rlbn5WORkBBgj13/AL88dzYh
aJ5eYqqbpGu8LUtEn981k2SAbEEOuljSd/X1OV7EteKNidCG1HzS+mWild0lv33MB31btx/J+bMr
Qw/VJQOmeCJQM2PAutdMYBf5GYVEXyui7LnNcNnENJyHRHm0wOzos+rUXKrQj+2nB7MJ/8i9ahcd
xuBA3wHmKLz3VmDmV5fIhEml+cp16B0IiSpGrjHyTk8bDK+iH647/0P29KOFcL0npQANua04cqoJ
x0Taj9eC22l88xdUQDjNUZ3VVpafSxrtrgQLpJbPXrA1elUqh3gScNWCHoUHeHycRofHeWV7Hp5x
wlUoHf3LODTtghuoA5nXcTtzqI0+p1rquCl4L00MblFoAjQ6SCAXNVdwVJ39Pdy9PAYu6K7nCmX3
OZGYwTDHzSmLVDJMxw8vu8kIsUX3fZqgeEmgP1CP5RouMkVSgPwlgKAhKoqfFEqJTPrfs6w2mEFK
p5qGvNDStKGEZVFQLwZ0EmqjXKRvKR5c35NVzKwZmdsxdoeoZ0ycr+Mve6NzZFHmpVbEFmGiZz+F
NK8606LE6OjgDZSw1Rs8QJ7MgHXsKC9ptIR4mMUScfkS+dpYBMFzJG414eOd0pbRRSIxyqWlzuks
8p0BkdWtAbP30p9jNPBzyHJNO0H08BlIuZrC1zTsgmMti2UKON3tG8YH2NuYA/NGWaGpSwQ124sx
/7AograCq+AwMBiO4b39272GsjxkkV+yenzF/uKGmVHPXZ7PbE7qCaIoTySAm3bzy+56bz7qejy8
vwWgc6qqRDceHzcHcLHorVxg7cKahraiI0dmjuT0UQXdp91eSV7RonhZnJHTL2pyWqPSY7eEOyv2
Wi5xk6f6H3soNrqsvDjiMhUdkYUzVRzwUh2HE0TlGHoGhVAqRShFexWmkltDhw4oXsWVZHunOk6X
0pOCn/1k4VsPgc3eM74POb+viWm4dy+TbPXM03FPGMGW/TWcI8lJ7UbcjEiEuCyf/SEDoT442LR4
4Dlk0amMqI3V6ag92tX5Z8WCC+wDaRt0PZqnr+prAYpuHgPdYf6WFmMskXzYE0yU3MBXmCFN1eqL
HQv+9rKrziaI4c3wYELjdbTtCqRg7f3Ub3/d8kUg5oW70s/6ktUh5gG6hhHE8RePMPCyNzOYezcC
gXLQF6G5ualwqcJlXaf/0MflxWNPInaPJUXlN6RCvHxedaCYT/pX1FZ6GXToVYEy4s2mK5xmTFcC
LfzO2s7i/r2WFvVs5NtwZoYmJskxZ0J9wk5F7eMz0zXBBxO9A6m8Cf/v9CnO6x+yYt2tyc4JeVNi
nbMQXISJaqfBw6mNIUGZXzERTanAH/riWrwi+zN8LYq3y5o6znnrfYhOjBd/lHydROLqMX2z3o7Q
HmhIooaAy2x9wy9KlcPZTUcvpKqM0bLKxdHwkPnUlsaPfmujbiFG6cBrXa3BU36aXJ87xon0xYsR
+CeGmZ/lAfB/7HD/kJokrUA4nNA+4ZTdlrGj+WrvUQoselEdUKZx1kinRJFT7D10Gd/Dk0Qzyt7T
/D4+fyuaNwPTpzmVJLSTuS9jZ1BIs78+4thFfX7Cx9r+atG+z6HFBnetYZFo0Q4xra0R7E7h/kca
feyfQa3wPrxWxxt/YWYIRS3GGEW8ZZvX4PC5lh0qkddYNju+CnvPK6TtPj+GrWA1B52xJdU7v0EL
9uHWUcKs/czTkLLq47Kex9W0SIMrDSsB7vz1/atX0RDCxT35VfMObbZNpJ/VyjzHZDVOTNqgcRYg
friit1Tx1wex2R7MPNIM9Ia4pn6GXWBTTOpYvXYYaq4ZyjVZ0nAZL5Df2TxyFgFl4FVsj7jkDe5e
Jns0vPCzI/xUIv2Q8WV7ck2LayKOPJwSyKB1OpsJMmfIszR5od+6ASY3eZiJFMsa1IPzzuKGvRij
OpgoP/SBMzn9D4WF2bPP3QZ1fZ9CVR19FbniPuN8fZyusRYZaEvznvEAkASj6An7bHpaSj8/T80J
97Z1bKzBuYi3AL010xiyxGUzpNwnyI6Oqx60c3NxEkbIhzbudyi5yDAm94VapXsWHXGXFOVmXQ5w
oIHntOMU/p/Ao+7sXb3FrLFIG8lhvnjWNyYyu+YiOA3h9pzKTilIJTAoOesadzhtqbI3+OQAyjYm
f5ioD+q0JhGB5pppFJmgHzzCZ6uN8Ylzdf15N1a/WEaKmn0gJMM5Ch1aKdcnzeXHO1iK9mSE3jtA
V2AmhVtE2ZcTE7ZDrei6YR3k4z2uz4FPDI2LNf6SinVENtIwlPyrOxDZZLCnYzta72n7c6LNLtLa
tt6isUhh0+DWcsQhKs5P+q0LuglBYZrcI7EaKY6IYvhopkNPvwGvEdp4c73TBocqXaqJMwKnAsGZ
6IieC3IyeOVz9W80J98Ik5pQId2rdwA6Yv59gh5LAM/KLfOwhqnAc/79jWQB9l9CtlBYdqwqHF1y
qULheeA5AGXesXrlk8AIj1HJA9uT6DN4yMjxQQ9Fhawx74PK13mFkci+zrAIdo5scKUmgHTXf56H
zKXHCDVoNhPhp6CGtnqnlDSW0XeqgZIl4VW6fqbTtvQqph2oFeODzO4KgO+zI+mdrsm0Ej8k7jKM
FK+TuKARUYg6nDebBulBVPEeRtcapKr8iE0gQc67zlcnAKoFmihC0q6Qzcn/9/v8JyvX4qbwvJkO
1tWzLyAJBACkivO8YIXPbscwAI+D8YPDN+EAMG7woW09PVvUV4po5/NsdMjFEWqJsvTJjQf8dIK9
qaILvBYBH277ndL7ZP0RwmFEK0Tq8U5DU8oJpGciTFIfhn8WZ9iIqfor0fBiaegXbsqJ/LZ94y8N
rbd0y8RYhEvJA3DpDwp80vI3AuFgYgrMuc7OKG+dGi1/5pSKNNZz7HswwoVdL/4yP5DqCeWt7D3U
STL/8l0hyC3uf4DQyUasv1++16yHHwQHqp9+ZvIdP9i2TvfDJ7SCDDz5KJJd0iVHAHqRIcW1+qYh
6SRh1iZx0e2k7jQmE/wS9vlm6yL3Rf1L2GzsS3ErctzI4RdH9Lr80XdeYG+qtCiOVm8V5BXEPAWM
gRxBFAlgta89Fii88a6g+tA8hB/j4mF894RuR5qBBG1GhNURbG8/jllGUmw59uoTkp5wKXqC4vXY
34glnZoPtIEb80tjteHCLFJhamRwpdFAb/+h1Ik0+Gq9r89zxK8We99sgV+++MCrG/CpthZtIknf
pusVg7W30nMgp1S0AyppdvlSInlo1RsnBIC9/cV7l7rffnVsdRgmMz953SAFMP2lVJItCdbz6s7i
wrIBZGB5WW5M7aEpbqLqdzZcdg4lG+IgR4wSbkzQDcafsmBxI5f3xg+5v434T1EmoHLhQDWHCNZg
9Tos3XF26xtwKvi/D+DgeRQeOfUnQTCyslzXfVa1HSDMsIHacz6v3vQQ9ExoiqIbPNqKnZv87+wi
NMVK1069y1xEPdCCYXIeXVHmB1tka1WiVWhaH8zxpcs68ureQutxz0Vs6qdKygYHrX953WZXi31U
ktBJe4ibT6Pskb9L04PBvh5oFfjgHne3vhJVlhCRQwBpLyqvPFzjsRvGDTXSdA/lr/xqfOyYqfKB
TYJXscTgzNL3MfOw28xCs1Gq8+X9kVWlTXR+NnWX4ldiVjim6awIhcR34sZuIeIE5jZDcmc0BQME
jWqV8xezXUxvkX59rJ2Oq166himsuNBMdbLzIRStKrMh2nU6v0G0NJrol/cClgk2onXGI8UtxJ6A
EH4qd6H2zKzHImDiYCRULVjahO/A7ETuwDtlRgnCzSvkBMe6enOL2EgghM+8FHrvNrjNWMzbK+WV
aitBakbgN6P7BlXf+gdfMiv5UsoV1pOrBvei26xQCUSTUgGYHf6nExEy52olSXGHVAkn7m6lBPZL
OH/Y+2TqCP5mpje4A1eo5F2gMD0OJbhnHTUnK+HRF0Qv2JVqqUxRQKhrKQCOqqrMOcnBW0MTj57F
iOK5oAOFnUKYlVrEJRG+f4W6WahKUMPHcvsBD5ng2ETL1P3WvqXqoXsl89BsGJWfAaVhPQFPOPCl
kSQqFY5xY7VG4vRNzElj7KZd1gvogX+8nsVa6IyKYOHVmaXbijXcfzak2YyLo+lDQ3nFGzTgOkWp
wlfonQhlQ1bWwhbKYnIpeaWRPVgWx0liLhrTD9V2YbsFXSgPUGJe6NGfzTJEfBt2wYaPXWhIetxn
k7FUHEm71sb9AWmmtWdwuJ74g9EBKLeM/gzIhO9ODI7M6O8dzS1BfzwSLcGjE/0JADLM/McvIlfn
D5QFL8HEayncIIL8njxRmKHYkoOH6JTuStb+ZsM3KBUbkAYu8iJLIy5ERZFJqay/BIQ5JVF381dH
zpqbw2l+Pa6XgIYQrWyVJ8q9FN77wVm3lnMg5iDQUxXujPBDQ6e1TOsr6I9lGBvrUYa/wPHXPeJ4
P1ufELMUj0ZGgvwqKV2niYZQNFHAJIxDOEN+vyfmQzkzNfmFnUFcEiYGP8i6y1tGXdFOGDbjOBr1
YSrtbd/UCFi/QlC+XHvMZ7dUh2cZY+HT+jYvwpoyvltLIAkxoYeXog1G4ho0QCEhQJodiQRBDBO/
zcdds8Zw2bJXISrU5u792Cdh72L4AMqT5C/oB+XpYKZIgqoeqIscVp5BbHghRKW7e+HD4n3bzV/Z
A8DVRxQw/x48AixzInLs7sYLEMFM0m2Yxbg6C3fZB1+CfVpwgDAMgP5oDuX/ZQfnbVm0xjx4sBdz
i6VZwzTdB/2CgyY8kDPVpszGkJpAt7PPCsEbPL6pHZR4bYgYDGkgnwauPtDpSCY7AZ+EqphHtDFe
I/tPhSISwrM7nmRtBPVcxnfi4+rqnsaPjzOhc+LcVXKVEwNrg4Kz68xPDyJT1O0vWcdjDWrnVshK
lGTWSEAwNbpoglbIs6CFW0tSM/Lf0x/oDXGpJm79AK6M+C2rpm+Xrwjt0aPrJv7wNa8JsAfR+Ixs
Owa2SgLcznhQjknX6ffOW5vW9u1kzXCMn7SfOyycKCRwyWtU4IARvHvyIgg1w5O17P5XWpYYURre
eC+iWX30de1A2VPL06khcTfuUYF/cVdtZa9trl8/77yIMpPRzwhUlVL92l0GG8i+ptEdNeavIr5N
KOKskYE5MzfdceB/NfuT9Olhyz4NnPjind827bGnTWw5/vCTEWkGmu9Ikyeg6rG76o2POPPNlMpk
1SyERV+x7t8KEeghbqsiuF0yfbptSAmJ81Gt1Fn8cxWNz1mCvse9Sxcs5CofBHZjWa0e7NT1Ewre
5VExDixmyV9ChWSjvNNFY0COa4BRPpcz4dpJeEGysr7V4a5W6GtaVv2XP4aFOeWh2iN6E7VHBwLo
l+TA1hCX91wWpZZO5N5ECKctTNXIzhC4a3xpPJA5biYMGEZlmPH/j/nwdTGKDvyDyvjukdb+VwgA
4hxFsxX3Lk5B2GYG0wp+x+0tJC38Ib4WxxBnKcnsIoOc40pDDPEmN+95oVedKcOemPvTN37eEDgw
w5PIe4Ch+JXNokdRZ4VwYskTDK8ViL1gTiAPcxxDK1TqpyEECQTtIwlT/+U+UAZVW3GEhAgfyVAh
KyGMdCnLE3msk7/+3JNBOTlzIWI0beLkk6L1a1sENpTPLSxnBpv/6ILDV3nZQfHiG0BemAlp78Nb
z+dsCRoZG+H1Xoc77a3qqmOpVun9s5qn50gUHQjKnTkRy9H0vkTyvtlrfClQ4HXzpLxVsCgp88oA
tmgdW/+t/bxRql72dVrZzTrqBkLRfVo4zu5FRyfN/h9dCohrShVqITP5FaABuux7VyCJISc8yfCP
a5rSDSqAowf4bU0UTnNrk+gDdSLFTwu2JZsIlhWpj37SIIZ/46FzC7gLtxN6D3ktfaDTYiNYkU7/
uqiuY7KYg497eToJ/tYE/OD0exUQVmJuYjLijP4svcmBoPQqJQL2uF8e7dnENJ/84TmCHAjXeTED
TNy+c48LBDMmmplJqnmFTexsGevVJyhsgrC25U1omxkE8vaRWoR91Y0ZfuAhskwHWoH6mGnSuAl6
mODP0dCdVZWKqn3Sm5C4jnpI6aPgU37ndCcRBF+I9di+hr6BQY/TwE/iFi8B9myZkOq5dcXPPWcJ
q9QB/PTowmVr4qeOtZ0sfMoEMQvGM6fPIkATFFSpuieJ6240mUetOXGkPj04/BC23JP7/wEzwBp8
hkrlgxQBWHQnbpLV47DK4xhY5hHZLlfbSaQTxQ/CW/CnlYDrJH6KHhKz4WeQgKgoiSWeaaA5+sZs
nyjeEvJzN55/6H06xRwwXCX2Fz7xg0x0XGijPMB4cnw+EdmpJzQ0QKwWylEUu+J8TSAB1ES6VDT3
zSi/YTT93mhl7k4bZif0TvY/X9g/VMLaxQ806tlU38Wg/eu0KtpyQQ7buTXB5RW8g/19Q9LZJ2IL
bdTGu/H4f6jJaZ3Xf1Q04lvMddbQcPbSRkF7zQAZ5QdPdMTTFZG2wS/p4QdNY8jF3v+HmGN8s+QC
3mCpEzASyB3WGeiU+ATxmytafBgOyLiAgxpfCKJMA2+Hwv8kPV4ic0FRpjW7XOjb9PyG9y+woyAv
q/QrigChacesVZAINHmokaIQ3J4lH6leucX0a5Nyeps/80Nbpa9rJPeGeVrS3gop3rup/KXn9z0c
w7TcA3WpcAM0/JAk9PAlurnFkFlOmenpK97uvCbjyt4A69R/bEKndMKLFB9H6ghIAAu+wWhRLaas
JJFmBmzVSrw8O8rCuK9jyTfh+g2btqLgm06ouokr6R0dlYVaiZQVISUf//qUzRsS7pKiBSBQUm8s
e3Bjg3Kk56RI/uY2uahV3ET+wg582IPr2KiA4ZdtrBtugv0JYVyqDjX6h4HpBNZtsRF1j1qbXxTJ
/HC0f+OC2198y1Blq1lehfRjbiSwCPF/+4mqCkBkznNEKENPKzVOuLX06cni8d+NERuwXb6fqRnm
JqUVnltJGIHUmMDVWqutvvcVICc3DiM9apnkk0gyrhDmudBcgJA9vLxeTs2g//n+/a1UQdWs/hfg
6v7atoQn0pkJKlfJEaNLwV+SY20EIVWDbQUqRXhnlveVdYmnLsj/hcqmZBIkva02tYmpjs0aY37y
a0vjHE9PSY435dGEIsfS5x89tQ7TaG0PQJ2CEgxX9C7xwM7MVX4tgAwwfOLKOfqy2N1MbyWwJTtE
KZB//9hlyK3k0bQXmXyeIVI4fzhA6bkolNXsurC5N3ZfYt5iEZak298/vexx+T+gsHhNe6cz8LJl
Xf0R34V8O74XzNd0fZOWpvgFCjUuHFtHnlpZPShu4R9GKFIDJcNTiaRJCtQSi6WbQZgVgIfdVuKv
qMihbRsP4Ci+Z+XZ6KrjKUVudoU7dlmrAvKWTIjNP0BCeRSwNVxDnibNgxRHs1mCGv7xDh1mKAB6
WdllcAgDCQWyBSkj57fBnPcqifGJ//NxMZSxNGL/zPiDxZNDwgTV8GcNLyJjhhqo7dLjZtvmfgVK
XdXJFsHWS9+tCnuOo465yCDtl92G4y8AwqVF39sJ1gt/Q6KwWTFcFZWFLHnQtNHUPCg2YYmvOkeq
N/jgdbeT13PNUYacO5Fkm4luaZv8aGETsZ2LQ1Fwu/66jlbRjJwIbyZTyJhvHv1PNG5EqVZ4vl97
Y68mQ8grfm16BkhdhdHwB4Ep8vG2tdnZ1vdiyniepSVpqng14WQw8sKUls1+aOqa8DrXlhkXvZAK
WR7IxRt1Pxiu3QS152SDIIqpERKYALNuhO2gw3ebDSOMzmrP/Q/pMoqBYaFvNQCyEZgNXJ80+hxd
VANFKyXL1UJ2JyvTzmnx8k+v+Q21Aks5rkLSMORs6U0fX1aj1GHPdu9a5CA2Or4zadktp/1mO009
ZjKUH9ovKJML2oM+Vvg91AEZn1V5nYOVz/HN/KA8b101DOxSXhYw7lBCCCgscKRYG3ZF6sRytB2t
k6xRDJgmHhl1Vw289yoXRRDfBOOI1Cad1XyNNe0exQEzv+s1Z1Rlkie4WY5tfUHGAAqAiPfAkFbT
7Ve6Dol9wzMfLjmeJ6tRTeqQxRsoW6bUyf15ekNQfBnNVSbU3YMNPpaMUKb3FGhUIHQ2o62ErLTE
8y5+PmjGPCdL51Wmar/HIVdwY7HGJBxfI1yV8kBAJkeOyk8lM9nuxXjYucpusMq0JTMKfYZ3txVq
bDYGAOpdcDHitx5GMKXQKKfkuynsipmxjEgeYknAeWPCqyIXrveLQzz1ninhaII7Wn1CXeoWhYEa
eV+Cf5epiuqj8CLf4AQSIqCxA7hq80M/nn7xoAVPOtdgLy8/Gckw/iE2K9cbMry0ng64y0x9DGRh
kXVInBXhckfOPOCH/AHad13PL/aNmwH74/2fN6z1fFOUL1LJF0SWwtbkf6ik3OjsiO/cq2I0gg2C
u+4wYWfEr0QAPdSXldgfd17SZrUA+xOpjGpio9YGeWw55IyhCB1vYDh1LBGmPaHs5w3+hFUTbp6/
khYD6oYZ9p0G/azdkgYbJKzJeqfUwI82d9PqN7uKwsFxu9xe9cb5mgtyaAYQElE8zw2X2IM1xEh0
AcD0c7MMPBk+TuJHQkaN9Rnftrw/aqei5fWym4b39vhJh8j2jNlfgIMf8SOVnlire+byKHkWwzRV
r7RLNtnYfJY9ejCc8v/932qYMp4tDeFPh6286qKwOWmrpEW/jgUb+aGOzMTwW3bw8BlY053hPGkB
sFmcmVnZpHCUyPLQ+hTikUcrBtCl8EcaDWLKJNZ4NMpBbNy/kAKzbg9lfUzitGyTc9VA23fapU3m
/5cBPLu8NOhrK37ys/JL2GBh9235thyed13J9/cPRUo6tkP/+fj33O+PPnrMkcDdPpZDO79zWEMC
FH2sTjZYA7hPpmsw3zHwHarX1inVXN3l0fQ6qwbhwuwFcAITZ7uJZyofPrtDO4aL9mD8XsHeq4W7
OL4EQX8MtpV2bn2y/hZNWgWTKg7smF7AzowMkxQln4QxEp/VUWphruE1z4wtJibVR8RARJxgPEg9
0k/a8wPU1ny6fpuPulkkBumK0deoEn9gsoDrj60jJeXIiUDPo5H0mtBWcZVjAqdtHmInqka8Ccpq
9k5wAWG5x6PXznNMzPoG5BdCaFbzb/oUW+YBgHK/zqbtD4SSvCioPsKOvcKejhTWwvpMXcufWzRr
BguqowNRxRds82UMvbswxMZF7sEjJJgL7IjXgIVmq7osl5lyVFIgRdV0vcPTnhQ6cyboC6L7/58g
ZrFnu6A8vwko3hz7t/d9i2wkBdbDHSaSFDg5Bq/k9LgEnbRbRVCtGrm85KjbhOO3p3mJrcBdYBQ1
YspXrfra/9k3we0deyWJqHzs1kQGDI3G4Urg8smTmnFzYZ7ATmA8Sqp9oi93Ure4JHS64TX8kLCQ
jPCUOTrNwuMyFAQ8Cb6EvTlopHwVC+NwCvOZMOi7wx/1KO7sD7xtTpd7I3bkZliEtrgAy3myqBBD
SSvIDqBUdgOySSTHuTIgzfRfN1lRe3Zl2sU2Z1+JqOO+bnaLUKWs0pGRw9ZZC+2aWCxiipOxyIzc
pe6CeVPX1n7jLrL7KcWeTuPj6+JNWNWTfyN5J9rhZ0owhXeRyDvwrtDDElNBYE961g98RlWlcmwb
6edm8PXYanOoezXHcis/Av5UUCn9Xb4/MIk34gCoV0LD96C7gjacKlK97NjiVBLwjzNYViUIDDFV
A0RYgJ2TIIF2imZ4YP4aDk77pPyczak84MKVhjGnjZni0D/ECKECfVBcu7JSxuACqqGvIIMLeUTQ
GIWS438Y3hRDF6wcvHOlUi/rdJe++wYm9KoWhz9a5JTJNhhq4BHIz3PNJTRCWios+HqOFGGtoOxk
8RZfjV0cPKkOFJHVB2b1thRy/p3NrM+kHDdYYbpfuz8X92NQVICfVkxFYBC2l/cSwfWDAglGN90A
zwJWdjq1LMgn2a1l98bWdT8uiLiSE2A7LtR80Zl7QUZge+t2Sa7KBw+tJaZk2y3OB/csd+vQ4+Ye
cHsXPlxVwf/TDdb+0PBJ9knsPM52eT8eAPYS6lCrAoMIGBQN4yte+gsmj/On4GGjbVTMtXlKYzVm
mwyeJqfsuaAyYQBNnbLVdVSbEiEXtpFLVl4sSaymtIE58qj86e1ErjUGDTW6msvn4sL6uK6q+zfo
nO2bHaEHQsFTcnwohiR75iufeiTg382lIy7qfFduNaIGH+dHf+ILAri4tC7xWFuMV28TItSkrCaU
yNE1PE7O9affHQWnlYkStBU9bcyGYWqaBl13+xqm4NCC2Z0HEQRnvS5H358HQKEmRuwvOCHw4o71
IrwNJ+B4Q1pGyYB6GwkojX4AO1q0fZlH6fDTPeTS8na6CfmuGs/1VJs4d5Zukpm4XiYFRZ/uAQg6
vPpFOdP8VNsuo29BExV3/or8TNBPBRK5D/dZ0lz4b+zNAzlZnJ7ycY6q009Rch8ue/CxUbOZTVVD
wOIS0Dmw78aAvNUI0BhYcPjMxm7UU236NP9bFSds0Kud3wfJwJS2IDLuMZcViBmL5qN+HSWBDAzg
K/FC5goS95kgVL35p1eDi1YbzHxlgUaeAtfLAsHbM5hsKyDwQtJcWOQQUFUesg7JGMubIdf0guTO
eTsXH3HqTuSNLNNpNjbfstw6TqbWJD0ofQ9oUvqovDxdvcWy34LrrMQdwFpLH0BS3tN/OjW3VcYx
rQ5zefbXxBX/H2r5OnbSN3YxxEXvSeYeNOTmR0Ja22hdn2z/fU8hosLBltS7dqza6md1RhCTUwaL
dk6SU/4wTYMNNNa20tyAlwQzxMsdvLELkg+P85HGimxVg8s56WnMKoIBj2cIqdb0OYDdh0V3MoW3
CcKdLF533Ycbsx87dSQrm5lr44XZNThG4ngAhkKMfFlhoHLRqZRR0DgOMFRDpdHEvR7c7u8k6czO
l+q3Wm51bRErya0CioCErkWfKNdMEQOZf4XEWwaPUvSFGW46DueFFJqGxp5QXEanj23eVCHgBznr
Nw6/wmn0eNZz5NiQK9gm62vKBew/A1H7GG+Xzq5ZeKoF5yE6wLu2VMzeDvwfXmnDV5FjVkiHJ4OI
S4qZ2djavHpTHnkONtbwhIt/8X79SZZj8PfagfYYpH5vRP3x5Uxr9k32HyG087XCpVB1iqZPP4pt
3jPDdfzkTmNxgxb0qRZ6qYfJpBNPv0a+wwdTmxSySr10bdv2Ro4cj13UQPF22+0HPynRjGwmXoQw
3uIhJZA22ygtqxt9H5m3u15GLXMyDZZDdTkXDYudQY0rlMsRnhhLgoWtcSUHQQs0boXk56GWXhdN
zjBJ2j6vrFP+c1Ugrje3JeeAtrsCNZPqI15hQoDRWbnxzkCs+95tqtpWh27XL3yQ+FB1YY+/zMUb
tv1yv/tW4mjHZ8lXA2TWZV3G0/AgDyuq2QS/+QeWQMwCLGei6ZNo827zDkVYGVPuAMKjGB9JOHUW
bCs1XmyyXtnOyBM0lbBLBGxHtxJYqWS4vm2f2fXlkDPzw2zPD2YX/89ISo0sOHpykfNt/1Qs0oIt
UHfCtilBqeLRe/kRcg9EJ9rEEqJdefOyLaNRKASsi23n+gvTWtJnimi6nFCE6fBkQyjlP+GH6sIM
nxyp/x3v91ViqU3Y8mWfZyfq4UDdC4yCVnLb7S1DuRxDCFgcQk0KWMzMJ5BNvWiXdRPXNg4Eu2Tf
ZRZYxKRCZxSnlTYw3IIBMdPfyvHFHhEhqeMnjz8ykLjxMA6142BTKRHRmUJf3PyAe6Q5mp5GOpT6
ldDgf2GcUdaTTzzszAaTvDYEc4Iu4JFhCpB9R0MZNYYk6NOzZp0xIOZ6F/9kz7DoyAVHSXmkntS0
Q4NE/Z/rg+S9pGLpVidALpw63jUS8fCAzj9Uq8FSQzcd+GshKxxm865cTBZCNM/qENRNf0bjOwDP
YlD7kFxG6QBntAMzb5m6rcbSHCUsEEZKMjxGuYnHJHdmVawlEYLTlajuR54+TCPdQad5igdMolcp
vxuwiZ/GZO10SF2U77vkkWqSKmDP6eZ9jpzp4UPGm8dBVj5dYxaGdpY0u1v/slz6aL/Ji38IgQKo
Hqb6mv9JoT0oEm+1RjHgZOX0+dVe+gbAVHRx04Cpds23mI6X8SW37mb5hHnRSlqpWYh8hT0ZdSK5
Dzqu5uPvg4FNF8enoPdW0lqA4RyqvgCqK/xBJ1rDSQ++CjO3e5K2EGgfjzPVKzBV3VVWGMXyDG3d
97T4MLSHRpJ/AfyIgp9W4N4sHYnk40FLJ0YEyM2l55+DNCSPmz5FUl6f1VGf7aLTC5txo3/ttmKW
9hAwf1df70PRTG59a6VwpEIpOkSVTxVbyTd+qMWANOmKwbx3rqsc0Qq13J3RqwF4LpU5MVhgxOD9
02Ltd4nwu5wosG+ZoxR70UuwQfG81/yaypuBB5Nv3doetdIFQTGjxq6iyqC+DbDtftIVpOjzkuyq
nW+hLcBCngTroJGMNHnNJjILxpkOLd5ngUwsmMVjpVVL2GNfC87wQ8MbSxj8+Unuj+ucnmSmA8dp
JuQfQpopeIl+6yJCIChf8C8Kpq75LNWpH+Prk8QxF1LCAOr3F+N4JLgPvnpewzw24RSturD5eI/R
TgRVldSxRXZFdT8sVp1aEBeXTGFU6mwlvpwzv8Z1aIMW3p8o9nDVxHNbdefxXpMeq1FFQq3afznW
qEcKHqt3Y/sxGlj5Di1Vf1yEXENDrUUPDLqYT1LttrM+SDaMBr45xKceNVy3s/T3/WOpB/ISGVdK
6qI1VEQMsAqzLqbyp2CK6kM9xyl9cWRRD4P+YY8U+rx2xuAku5ikxvwdq/bpzNCOZrjxfeojNGOL
WitMlj/sp0IGArUBztFpymsbCpI+gPtK2MYYEFnXUWf2ZuCaICHQS9HK/kDbHxZ5OH4uR2P+MkRS
X1XfO4lvia7Ol35VDGTdr05tV4KyUxBhafAa7dgJcWDkDQca8TpYBzFZeobGJ1T/c4/+zhIpkE10
BX5ggJingIDDuFPuzzr4QfPOVAditVcpkfHFhs6aQVhKSfizrqmxkt5q62ytBFOT3wjLqarBrDca
g81jghdPo2Kyl4d3PmFKag0HFEj/yYkTOdrdxM4o0I1CfqWZxfRoN/vFI5mP+nCPNoPrHJtKwXpQ
WAKHRtyYBzjUhs/foI1NNas/AfTpLrN+tiXUjKt0qfkUSaHfAaU9HwPhwPQpc5mjGXVBCGWEQU7w
/nkTCDuiMMezeKgt5eUmHOI4Fi96wP8FTEoB00RM0GT04OETsAPIjEu77waOy8P7JzwbA0h79oNO
i8jnvi/5Sj4WwZiDI86KUrF7yCZJX4nI65dR053TJ49UR41G+l4MadH2TvJFYhL1+HQ3yJnN0ptg
xvoDBFJw4fRwo5rw4tj1iPY5N+CdXBVy0aeHoglhtlDhB6qOSsz02Hv7xgbxnYFGPCmvHotrO6jJ
NZy2kfvWbQ9Byw1xO3O5q+OqFO4xCEuvx5eC0sSUbLW3Img8yiPY+LQKuPLi/Bpz8sC4HaTkoLZO
4DhEmCf7gHhCV/nLQlRL/EPRvygV6cdp4RTmdnzXqIOIDjpqTSP0Q4Rivi4GcNX25h+MHmcw2Orj
5s/RIPwmza+Z8jUI1zhg57KggKHsyX0M+DOKj27CAivFPH5iZRzkcmnSc4rV49DSAxEY4+qFbOnR
smngWupWZ72gqJuDbRIX/NUSgrzyV/5DB4QJmrHnFRnsa978w+eYFzUbHiBYtjZCPehRA4T0waJU
j6uX/kaEXhMBLQUmXkNwxn8qjp0xSfACvjWKwEelT/Ibw/n1OrQgK1FoR26TobCIkTEYsXUbftl0
GoCtWs4tLwDTsc+fr6keZ7RFjfpgIE0cId1FS5F7XeYiygEoQW0iUtYT+POnqYJuHdLgA9ZNdpEU
9GVFbuUhBrjZg2B9S4QBEFuhKQmCVm2QHMBWvNqcNfyGCS2kLjtf91McoWkrIBUlTbRSyhXsz0I6
dPuxmbfvaiN5qCGnRldls2qsbgWBxB5MeoGutb38Wc3wKMmW/+A3ljfkHbk4dqFjUV+DY8VrssIb
0fnN0Xz7q+wwoYCSkW7+TgJxVcMV/Y6p6eC5c/+wOYofy80+eEogr/qJWEfNOld51Do5Y4MyYWmi
bj2GICQYuh5mLgLKbdJlwGlxVB088p5Ki9VW2QhFmJYDBtWPDo+5Gwd/ycVj5uKmyY/DwGlgrZRS
kJ3N/DPlWm+M4NDxoL8Q95O3E+tmWN2FwN06oz262n/Q5+5Y/yP05oxOQghc2MGbRL4EtFKq26OJ
2UaKUNaWSCa6GBCoovq5CL8OyvNywaGM2VZN6xm/rSA8EdFsyOfkfhK7FkNxalF4aTMLpBFBqXBn
iQkeLLewu657m4mJ9TjcYai83s98c9A0/6PX7esxlWLYSLIIR7HjR9yU+LfqBVmUEYQqYsBnmKV8
eHPeiGhwHOhYUM1SWSEmubS7iZjjvfHa6jKKF/3nvdXye0/A5A9+3lMKA9tA5b0BLhP2JuLDZOxe
+j6bacvuJh5ErkGLeJLhj82etAdIu+K9A5RYBFOfCg0KYVMw9vZ7dVytBgEZkOnAJxTj/S+UYWCW
jkYluiC9f0/nBphv+hE4fngf+OjVkrr6R2tcP0mFrmNMRuxHDVAtyVVE08BHSb32/UCG74eR6vyb
xO+bwjf5xu4xrCQhSfnyCTMwZD0HsfgF+XEQIFYeaIcqqbLWHVlLu9mJ7hkmfNv7fC5qoAIm05jX
DKlQLui9KFuuXO/yvwwsraNWLQpsY5jXlf98hhzC/u/DMmUd4zRkKIatHg6ow+aMByk8hSOCJFDI
YA2N+v22rRqPKGovp2OSvQDo7FwaZZZC0hmF4kfVT7U6BO/j/7l3rqARjkh98YkmmEfGTsp5/MZa
yp6e6L+2K5Wl0/jE9/G6iqzsJAsiD6oO17fiEjvJ5ZamzwiGWgN3mdQRLirJSQV5NZdUCBnQJTVq
7q3R6FxseO4W9q0Rs26sWlIQ6MbiXi3okAk60W6mUVjUqwLQXsJjjZwuewIGRM8jdglWPKKf4w14
q5HTuXcvbq02N+leWlZyzLlh2AmnsUJFYOoKqC7sRU3oUyfOU8lOwoWRkQV7l/8s3bEzWykV0aKZ
ldNhXdV60dedQ7Q59ULMofCCxtbHGBcUX3/8Tagd7fWgJWnvposAlykvNiYB+of/iIrZG8EPZIta
SE8E9yPJqZebd5G2A58bgKTh1+pNQSd7UAnAl+9WruOHpSpOP/+r71dvRsKgY3YGSYczECMtl7ip
lESE9oqPvX+5EpUHkykHRkP5ntAp8IxmI9UAty3VSNrW/x9kcakiPBe7uOfIksMVZV8YDr6FJ/IR
mA+e0tGT60rwsiFBfvonqeUBYg6rfFe+PJnE7O/ZfpSjG7BnlVdnrWa12HDuCzjQWkTOGFCTVpOt
6/Na0iYm0yYPGN5oYVXBYTN3MaKgYXZ6bJFhOKKguZrZJaIyeNjS42GgsAoy1r4Do2AkjhY/i6sO
MO3vUf+vccSRWiA/CYsBjrtXr2bapY6coEjb2SnG2otDpcKVR9qJpmUW+SfKb4u5V3vJp5iCVxP4
jBiH0a2E1DCDZW4CFIXCX4EaK/31Zzp75tKR/5wFQAORnOU63rdB3V2Cx85qZPYS7Dpn8TjqKxJ0
Y9getxO6Qh4oicCMd4e7k6nO5Wqg7czFNeV0cGPviw35UZBNOLSOL0pqGj7VVw6Rk8KywU3jd1ec
ak3RXZOtAVv9ylU8QL68cg/+oKBpMsA1IhXDIEP0+xK6DCoO8uTZI/rEbHQD54OlX7vhmiS0jLlm
+E/b9uVzptMZ889MqrAKLTw9By3qOibHqVGx8B6Bo/HaUi+ALrXK2DHBMTj3VK7D3wpALKjyquzF
PysWiXmwx+Fe0wI3lB5LAuWrPKRaJddbRzPZ08sKXXvYnD9Bz5EILxzxUYo7NSjIHJ0P++saMSiS
KfbkK6sf0Yr5ZWrPftk5MoxgIPcTAYmKcKjUX7FWrh04z8EEa6x1RRFJEt2gcYpll1AONBmeyN0E
74nbDNVPOcDzQo5ajiVYcUrCsXg8OXAI364t4NgfVFQT7zmZ4dlw5FJGXW0yKb7UMlRoh/Hkn0oG
YBYYvbYlcJjdpetJU2gji+tjc5fUJBmkYP8IuME/T+vrXJ1xthmRNHVBpxUKJrwbNDGLPCHq2O0j
v31SX07JDQpeR5TQBxi9ft3Tx7jQfoBPbE7Cy6gc7yH9D7jeGP1KsGnhvufv6dwZTDbjaAQfc3R7
gTdeXYba4jclxnZYOy1ir1kkSKA4DCU/yznvqaf1sJ0qI6qNpvKN3W9Sh49v+f4b/VfnN/mFOStS
m+vlEWpDrhQSgCSQmaf2z5qNJ5qaiclnZS2o+rh3jH2qEWhoH0do+Yp9hlADqFO9o7cYoGKJRzHw
8aUFSKiJ0MCqUvFvXISwXXhVoxBOhCKbG2Y6C3rctkOT9TRkVctnC1Lygq21sMgytRhAkbTrsmer
IOIg1BrE6QAqezLON0FqivBXfmayvXDpPSSIDUoiCe927+38dUm3fKMT+RauLFi1wzHmnNcE97eD
+X4zQKX2ZVjMO99PMNof4oqQFa5kesmz/DZEyO6Czwhfqb0pp34eiRSzHXB6A/Tc3TEc2lechZx/
1er4nVcedXQbysz/GmMECeUwPrxahtoTYsriupqlquHE6bXARZF2RAMsW+K6QIVeXbCX4YR2b4d/
R57/My01ZpyYyvfuoRdLdeKQl/d5C67AX9Fd+Z6sqeDojgCNqk50yzhTmsowEXLQ63chJ2rYdchX
p/PwNYORbmOOD9jfg2eLG4Snd79w4DI/ltUDnK4W+8vTYNatmouja5f1XRFEq101var7YLfSOjG8
jlTNNmhBImBXrhL7qN+kBlxq3ID8ETG0oUGlhHgTz7hF6N59L5UH7U1pv9e/ogmFmh/XkC6cenCb
71pe5zVRSi0qVu5Y/Rk/yIK6ed2ZyqAW17Lq591xkWwuU6rAnlIaL4rxvng/7DeNFtZu2lQ2Ha4p
PoUL4cGsiRHWKdcld69+BYqthtfuH3M2g1PC9gb5ETCkUm9RWU5IN3nKJFJbyQ206csglTIcwQFO
rCAelw6ZuloWwa3I29MzglyAOC7F0XQGV+2z45Zgfg5kJQSgF14aDWNoXCHQU57bz0sD2XpvE05z
mc0Qh3K8EMV7ZaCtJIl6KfCSHPh/cXIP9z+2lzSG+qeBAHhaUJZJJQPfjPRBVrdv69RmLD75VEW3
+JOWy4xo/jQDfdOyBMts1d7jpNXdZAayVj0YHf0TNC4c5SThpoR6TUEBwVUVwRjxO2uOQRoU/Qaf
sgwetQpN2gKhFG77dCm0VGMTrwnSqCQS/ESf5feWcyBK0xP3Ul24gJpFJUpXcMigB46U6Wvz2CaK
VpP1y8rNn605QO9gBLnWMA+sa1a5oLPSQGv9ptWkMMXRDz2khZfPQ14bCYqNzSx4rEhEc6O8a0W4
r10yhUnK4ZSbH/Aqu3LoAxnPk/JJ+3GjxsPP5uyDZ/jOWvOjBwyXuGuS4Loyy/BBQi2lAU876x4T
dCEDhzRXCIxRPJNeMMIIPTLztQpJGsB5L4B4ElAKMJ6MT5xMpery+pqCUzTJDWQvtWu+zao4ja23
5cqkR1qk+AHP8IDVlo6JmOMSJmc0sJaX5NrP+jhNxb4YdpDmWbrhkQUkrhyReme3hKsrzpOEbcWh
+SZI49fWppK8WQ6tEJkOfN6Z4ALMuxqv8VUaE+wt1tyyGX0s1IAz3JmyoQihKz+nZTV9hkoOE+Q9
sU2y4AOUMpmATLHPSR438TvIEMMNPJ5sCJZFOI3PIjyUZi4YNNdeczG9osb4UnMu+KC0knN4PtJ6
ZDn4cfC6OIW3SNtQWFWEWkNFfBtDRJbs9prx+ki4GpsdpAG1O4z/1n/tsuhiEpxH3R0pHR3ZBC3G
jd7JGWTdmP1O6ua7OBOQpybCLyEId7chiPpK+MauHLC+yxrjv74vr5rzYGz4ac/u0gR5Seor5uhW
tsjk9PAtgqtrzxFeZKbZqCcyt+ulGSPScBLXZitE0hnAgjQbHVa9xr369vGKYrLqeR4e1bUK7xEj
G71n+REfXfdO2EPmicyg7fo9mdxJkwQ4Y2w56+J2NncT7Nrp54I9kcljLCrggUJB/zSiRYcAZIOi
tVnGw+Bb7Bo6ekbvCxOyFwmRg+lMfzmSjowah3VZ57sRpNOPx0m7/73QrdUF+oJGXpJ00D67rf3D
G4Kyf6Xwl4egi92ukIEdA28fcI81WyPHIxfcnqoQ9gH0oIa1t6f/zuSx+1RaYx3cMNkHNwnNyupH
k6XckxtZOc3svY6iLgVcjtjYQ0h3Y2y281IFGuRUO2045L0Rwx6vxw3EMjQqBtQkVWLdAXILMNDG
4qAvX4d85rTXGAPl2KQoV0FYEUic+GvON0JS4sB6SmVg9OQSP3lr3w9sl01KUOgTy3M75GDr3jql
O30qTmO+43W5jQc82MNYyPUdx/mfKdl+73SVW4XeyaMv1EoLgj5CpDBv4jiW3rJO085bfuwOGXoP
fEc22nAqcfGhbVLzKqKAD4Dzir5Sy5DdUp+R5HeLC/qCEl31RVl9miG7Bqji5SMnnZDrkIWQ3YQV
fs2m5aLfy4thWkZE9tPRgXGCo2x7GoH55qHZmNOmJXPgg9ZrSv0Ko3Wl0FSNNfDV0M6mra7KCiUC
2J/g1IK7oqrLcE79q9iihcQgfApoquItE08Bj8rGS6HJ9dvBweyzedzEmpLezcn3CkaE+bRx5clc
/Sse4YYoNPTsaMKP/1P4A53I8AnIWkhSy76Y+4pGRNrkz+VA5GmNaaPQC+pZwVY6chlL8MSte1EX
ZDtPDIjjiO5nwFQBpoef/MTSUCrumB4zcTBOmuSdf9l1I4ZICX/u60DCNlz3cNL8dbi+kp39I4+h
x4Cw7J2MUiKt22cbH6r7/v0xnb5DlYeiklh8OHO9dUufdxzFutCyO0JbennrCi9MzjpSXSAuThie
a5++iDLsFwg+7TZhykQuj/Bv2SHm0vZFZad9GZ06I2g+rqzLp3wo6PaDHkn8P8AaEslTj76gH/JV
Jn2BraiZ9Rd7AbR2Ilg+y/t4lixYchTRXh2uynhRWICWyL870ApZKU5cmAVFTKK+CbRHC71IjWu3
AfugeqgpaxrRsWrgHCwaEyERIlHmzLnUenKX6tDc//c1Y66pGKJw+YtOKNNkWs+U7Ln0uKlfqQhb
+EBZYu4g8pYA7w6R6pBKe19BTvOKQm7di0K8Qe/gIW7tay2i17vyW0XEQbHjumX6Ifzfq+knft0g
YFrovGR1KYNr5b/ax6q6aUmV7NgMFUXItoMKbs9cTkwMbpWMv810E6y79teErKQQN4J+8PLq/B2f
aW3/UwDpZ4f+QD7FRprWYqRmw+BE69eMz2TZVCrAQ3Bd1O3FdIr5KQNMQyZuet3RlHlW8pzoqnOy
m6h3In0mb2M/vtJTud8u1JqK73pc7/9NWBbDZQIodKxmFVfPLlZaTn56+BrSZyEza8wNO8svNVP5
FfocIFTdR3oGZJLN+EurFUiRWTiP77LYvte+wTLviWnqv/mvNn/K8pCsTiIE47M4gowaRspybck/
wWqBvDyfNPD+xYgVonCmd1AAIe0Cc06bNPf1ChH9GMpVSCrp4GoZrZk8aLKGIcB8OnyB5H1D7YSp
BTHoycnuj+ShovD35SyEgJQhRSxgbS0BDMlKYdxU+CxXi8bWiqSSI6UceYUkTMLdc9aeNr2GSKOp
p0OZo/fB3l66myqEEaXqyxFfWnCHmHt50VG7xm6M9PDySsyoHeYe2ebZRpd25J3n5oCT0eFJ3ueb
0O0fU3PKtW3qof9SkgCB9njJj0P589xVRiLFUbR8u8Dhg30BxWjBt+znRInym5lsq8Pw43FVTa9l
6q7aeYU/Gz8pw6SwKikOdUcHf9n7ybJK3R8l4AOxMIO4Lek0Fj3ltW9HXQuJIy3NVub9oLvTk4HG
ZZcCZY6oeJH3M3vN0tdQfs+KuH7+HbDRX06W+30RqptJvS4syMG9sM9LYBitO2F2Yg6vrYDD312Z
y9PnBUND1/BxnQGRxhZTv1H3J3MBKu8TDTWivO7WFTYCA4kMZoK7f5IOu/q6Oe/uWg7Anqi8KgR2
SvJKfoKM/VIo9t9be8TkQ6V0cvZBFADpdM0RqeoKf/h7hWMVVuhCJC5hwsTlzaykF3JVC6zfmJLV
EFigYcXEU71v1ZXnFNREkxU7owOSRqRB+1LNJRx9zVUufGboaLr2/i2NcCItO91qyH/5a0oyFK+X
pAwigZA6XAeu/8b85JMg8dQFo6+GL0U9c/pLvVnQR7RgFtJxRjisgCYzxFxE+/goO3SsjkU5nirR
cCgV90EaWRPmKgmGNdqWEhEolBVDHAiYMnx4t32viWquvYvAIVvgmCtjp7R1Hucrf7VgNpk6dA82
HS7Lol7SErh+SOOjKzmtPSLaKii/NMdZbYym42CiD+XkRb+ECtOmMOoSqdVCz7frgKFDMCEAtP6w
N9KAHHBY5RmK8KEqRsGR50YPZ4GGEmCnEC08hlKdYcfX1h5NXZnOfM//L+gGTZsNlZza9fNfWMw/
e/Or/w/8C6RrAuz8kyzMk1aXLrMuV9NAX21NkmMjqQo7HAUB1Wa6B3jF43ptOg2PhksCcC1tSckf
CTV258AT12Lh9YfL/RRp3xS5cO0ws+uT7NjQeajkzQthROxApnPJG/Zlot5h6Y5/nksTmVScQ1Vd
h6CTJ8vDGkYv+poHL9xvm6xfxy6yW11iDEkzRcDjJJLotgNIQsAndq7SgA4Co9cKKFBrAogYDcRT
WgV0JuLd3wi6BrFAGoV/qHZdyasInIFQQrNM2S9crpGY5vWFs0AVWgiw4dAuPCMJ/a3lFXo7xBnB
0hg6hQRWHnnGenOchMFFM/q1hoQ53MHCV9gKEHZCrQXuwGyCffATORxAMEXMfgjwCjEa0f7WwwNT
UOZUpiY2co0jnLtmMHqb3dd8KewPZzXWaPTTM9nhDU5axuS6LasxxrRCH817XL0sjfk2mYrBPOY9
EtDtToIAOOT7H9lf8cwmTtxN9jgV3OH2yhBPXujj71Svg/7VqVlDf+VSoTaL2MBTqRrxhSORDlxC
j69MIP5psBb54cdGS1wt2V9Jpz9VI4nibI6EFdLsbkdNoVoXvPb80hWiEZtvzt6Ql2j7Hf97lMD4
RmWce0Kpqj7bN/yscMWsuhRIZHzc1+65qmdm9jV1hh69tzkQcBI/Tn+d+aTjWAffuEKYUKH/v/Ld
OAb0WgSsHKoWY3vtNXwNQfaPpRHxa2sgGxGW6HCZEyQnp+I+s96Q8qQVcxWND6FOmHm4Nr+hcyxl
/AUraZGzbPfIbgC6+iaDiU1c5ENydOFSeA1oUNwVeNtfiPuWt9uC2TOTOdr8I29Jq22lAvmmrVyB
IIU4KjbrVWe7Xr4lIsLgCK5UpytXZPTmbeJT+nT6AKmvyd3Lyr9o1jDQ37Vh8vzGfQvv/hIJDQib
U2e3c4wSP50u0kMTaKnV/g0/hDt6+HxVIiHXPuTnEiJDK3SzqeIZTNeUkKJdOGGYNwRAvrz4C450
yRSdSmBluu/p84L39CRFBUVb9ghJlGHSOfnhlejK+IArci5n/FlQGYAKL+xMd9nI84owsEYMx48w
eI+wSzhGomWpEZYWYW9M/dHo/DKULAIf+e4IGSoiV++Jbn+y1bTKx8LX+hKc4kwHwpSN/QZl8i+Q
fZn/WUWt4gYy+f3XxIb4LRM4yGhS2hz5yZyhXg+Rbqt7i1OpyRMfI01v6WzvLCAd4FsLQFgko1JL
R8RXz6HSQN+VzWWr6rJS+IZOoolVJ6Z6TGExxX9kjqM4yCGnSIdd4iMnPnnYEFQOFGaybhh5uJ4m
pgsdtORrQ5QDsbwKv2ICu0ZUv1b83bjAbkot8dA4tURPR4kr2iFKzxA8RGvDCckdp+PuR4/95wU5
RhD9CoAUP38hAnIIimvlCmJwqqPrw4FWIlyqLv+6Y3QXt0WIrgXSg8g5cEVXCPPpK626x8rufkQG
J/nJW0sNrzVchV4aFsvkwFaPkPsytwkpQA35rGng2yre5OAH3G2WDEWxl40x1Fl38qtQpRkFvth/
G5Agpz3J/iR/mT66tgaF93Y25aXfDnRcI7r8tZ5nBdvxS9eJXolNDVTD2E5ceodRCHGSr1zQhap+
fQQrGxkt1yvqZKKMV5aMyT1yfV9VAbhpG7UzPh3Mts25y1+f/whCzoDp6/os2B4iXZvH/cpYUCBf
dvv8fpzwYskNGNH63EWxH5MvC2c1cdvzBIcDEd4e30Q50uKwkjVqgY9sW7N8v6/luJ65bms3J+6z
UJwiuTdH8ezp7a77rUTsh/Oy6m0y/9hQBwCPuxYCZmnNiK6XLThqhqXmomnysaO3UYZHAh54P/G/
jGV6qVHCK6H8O6ryFoa7uzUYETFo2MngtThFQPcHQbp6u7dGp4GWBVP6GxYFmQqZjSB85VSdu2ei
kAIZd0r+z8SfHSKsOFKur39Ms3J/jkgMxTqhptIsRxpsAnlhDfEK6HvWjPMq5J/QFgX+hn3Xv1Dn
mwh+TXW9Q2Y4drqOrmB7F3tFw8LwkCNljvwMD4wDYlz99VSmqR3ebBhkyIpgJCwFPunJcGCTfZ1M
6zXk511h+4ePOfsYSlE8ha00SWKITZZKUxKuKqxuniX5KDTmWBtJpis8GRk7H4wUDxuPXLWq8OhV
MCeoiLOi7PwJDjje6QxK2XHnKDp5i9/dZkhVNnsk0hhdqsXrAwFF8oyuU+YlsjAtbFfDxujN8zQw
DEdl5yhzeSYjY61z/sCOe8fxW1tEbE6j3Crq0hOfWt6myhJ1uQRFAnLs7NxEkOal0rAMbHiOFh1Y
/99/a2XLe+WPFgaLZNL0YFbWly3jSMd6pLlAeO3Fvnex65D3UWudE7+6jYCkqyn8QJ/iLIZm1iHI
7vwDJBVIb6Ne9GUmTaOB1sfYSSO72QMLAVteYROPwZaHcXXwaJ8cxIbIMa+UCXV0LGmovFTPtiyc
W2StrPOZypioBmjZk/CtWZFGjcqaVZ5EpZfkS0/r629TvZ/AcRvNtkaJrv1CqcnuB1lKX4GWAMAt
SYKo/1q59dYkUi56m+D4bMuUD6S0DsmnwAj7Yc94bLriLrwgQ70lbWBu+H5OVSg+sI71nxtC+GzM
7E1jTw+jdnRJ5xV3eya993DERXvF0hOM7IakmoxReMohRYJ8kQKQi1nmbI0ghvziKJRWWhfgVfXO
cqDG8fQlPG3PX8jcq5w9NUWxVUTDcEwUkSPQ98e1U/aii/EUokLiIkEeOW8fJh1mtWH57iceYeCJ
IaGpnqSKZAZnbn5aYpsh5DWH5+hMXa+txtAIKzERoKXZr0ffHr6AREChCquYJw/or5Os8XChed7C
FcAuxNNxOaY1bf7EpOLrZfP/1+FlfIhbLcoiS2Yo75rD6j1tiIry5Asey6C4S+0q/6OCND2qNOQA
AxQ8KqpU/AMcCqRrzxSHk17g/hFEY+qp4pxNWofWJmKIc2bbSlfTM6l7V9rDQdWpxK5BZpHQi0yu
A3R0vKwUQ89HMPf0aaS/8Eb6ZezHzJIYsbArLKHqLMyM1wfty3lIF5WrnHUnO4u1Uw6HFuVwUKUl
gj12S4kNDap/KCwbM/EX01MUt69XzK8nhaCPlZVoaJEfhvjO3MVRtyse/2bZ9UNu23nUNm+FgKbb
rMUItkbbLYza/qCzg+GzJTzEw8euFOl6jTxurB1f5spnhGYfwX8B3bak0F+i5SDuhuc/Oo9WdDrT
peNdu1YdU1kAXw8rwkq4KzS8RQCAwW2YIIYyjCq+dQGiadvkejdfrpHRae6fHBZWF159M67Jemv1
HnApJ/0vwmBOW58XjQjtUh/NCeAZzVsrBeewZSYJsfXGXn3+AK1gRqFWiYz7+jBvHE6uVdFwhpM9
cm/smWn66zLH7rrdMdHym/NBGNz4CsWqEagB6pZ9wHAVskGkLAtR69fJXQs06T+n3WJAjCn3zbw+
gVz/T7d6am+VBm0KpoIMF0YZRpgyDxeiT97W4wzse5rnh8Kkwbc/yOdmcHeg+QVzmfdzYq+rauor
6DLkQmyYEs6Re6an5vQW1f1fxB1POBhiqRONrTPkebxjrpe7GEv7y9g9MA3Efp6feAjlsSrtPkYO
7X3ZH2wGrApUz83XCqYOes5D5gDzZG0is64h35ymkhZPJ/iLWouOBafrLyXU+0srj30BYHlAji6e
fWibkvUmMh/XIFuYqflrS+p4aobpGJhSbImV1lWoKgzH9R9fxvyM8jgEC6D5iG148xHa/q8/vzy4
9uU7IN5pUz+W3kdMnnCzDWjsnAKTJf+KgRzHK4EdSYE6XaExilV6zIL+RUzTpp/TQ3kX9EIaBupV
oCz4tk/+UvCJHyxsy4GDn0NYGRghQVfsfWMP/VaUUHw+k5OE84llz3VDkfHgU6Aj/twe/aV0L00L
9h+X+eA15R+BxF3ogBDLmchB9dbmaC1WExPXaS+DA3vhGDHs0BFnpr3a2AyCVBJ1Hi7Ws/69hSSP
/d3L0nMtIJpvgXYI4MO6HisHu4SDgWWCq9qhw6PDYhq68p5K/oib1Me+1dubAFthS0mSxC39kx6n
A0ym2rU0a/nSrdPpAj4Sq588GftcQNXDJsfLd9c95cDt9JCs8AsaBO42dVRQmiNMID9CEs9XTotg
/9b4y8TjVYzL2XJDUsWoR7hP11iqhRzpo+8Rf+S9FeUXFA0N0igJ8CviVl4Y8Rx/NrUXjrlgdJhZ
lUbtTLRsH0ye4ENzxBzGOcJNFEQNWmjMn6uYSshuF0hBR0eUHjpCyPeTXD1WvrR4L413BSxOgklg
6w8MwS83vOW4Xwwc2jX+ULWjMbtfyRFJwZ3+UQzdMk0zAyXhmqOXtWX1cap1wslzLrLzYnsVBj6n
0bx5wcW4X5TLV6zKMpUi8JUi4ZxfKH28UW6BZj91dPeDY3CriXWejdGfoeNJP9dPgjE2O+U1XViX
ILqvmjNGuyERFKSPcGAFXBmYBTc00dYY2IByAU+F+7loKx8sZfB1rRcGP1/OENqsd/P883uKyODO
oIUMYKwFQXo+fUraXmUQQumiKJR6hYx5gjbjw5pdTTzruDo3yhHKNJmqHzvIC6FxxQvyN0tDFGUC
Ck5FUMOv4uCXpzc+kpn03cy1d1Jl5AUUz9VTunZ+vWFabgez295iBis3yvQ2eEG/xES2t3vmSzi8
rF1/BB13019/e0qgxKB1ZOovFNyn4Hz1aIw0/z9sK1B0Z1UnsMUxfQb7qSLL47dGsiPnXI9Z8hyT
pZuqt1zWhgfdwv2HFBB87X4pEQcCMwfgYp2iACt3zhCc5IPgzGVwC0XkBoMxSRLWnakNjUpnm9JG
9nUr/woiAnE+Tif0bf/OmED6Mi7MPDX05aUsBptHHmu04u7VmEnvQvwGsxFsqAGyK63uWhn3zL81
ZtmMZMTN8n59L6xSYtmp3/8tUJ4Sy+m/xNnap+A2FijbcKYDCbwqgNp3ipqLX4Gn72ONQDV/PDAi
Wzgyo/GAw2rWkiAL8NXt4qcIrg6ZeoAaQiQrC+ih2tTjHGjrf8MrFiwGSfSFWigPLgVKZvlpANkL
tLPoQwXPae8o/cTW5v5S0MPXqkkv/CYnxMGSSDNQv5zUzhEifPx/jiEkqbaxt5Ji0Gis4pusFMKx
LTs4WWD7Zo3O5djTiv+YqVgxNQJ8vV0Dw/dPEcaLXSxoEN82qQucg+a39zrWHI/JZuQCpIGE8oSA
2Np1qGzQspMden2iaHS4/pu8I8eEEOa1e7WGXH7OUVOBMtjk2UDSn/GEe53Uhv2wrmjCQA4yMR1B
N3EhA/cmXIm8e+Yevk+PRzVxML9snxt79dya+s+2i90Pe5aG+G2mpTFTKgG5J2DO0C3t0HH4FPWH
u9gcxZNvGGgoNJZw+Ksjl17phYnnKJ/DNglheQvg7pxJbx7FS69JPUs7N7SA3XAZjk3/Ws8eDhct
XuGPNnTiKuUBJfiyl0deMsw9c9i37hR6JxZXXVXYEwmWcqoW01tS4IaL8aYbuVZ8qA6SfifOA43T
83NJr2j7OU+DsxWQB81O8Uh0rSJlvG2CbnMD97cngdREcp9q23IgJUBsbDlXvxIdR7VPrH+Tp5Gg
U8Q2HflutctI1i5EdYOhKwm/8kMkQPBownnkJdbRoSuqB8haEgczBSrv+Xgex3y2eKol/IGdu73O
VGP9LgWfGYR5icOLqbFW3fTqLBVCoRItZHz5ozthKFRC9GjKe+M1CYD2aRthsgOI62CFgTOsu2Cy
iBcFq2UpPb+svrYr6pI/bvZfQXW/pcwuPOT7Yl9333a5QwoAoZd0tXlZvSMrRIJ9BmcxBOqQty9u
Y/310eosUgMoMnhGVQOsyI54wDJz9+oHwh8ZB53SbWQCvjdqHb0XUaLuzpWCC2YHv294zQpuNSNN
Ixb9cBjoo83g9Tyupmg2dKAKySRMhUsW/hvda7J9JS9GCzSOlMhxCCzg7I+y1D72rebL204lbqGo
pDvp9JaTlqmXqOhF30HASEsF5LradtnIyqbkmldiBPx8vTb/h6igufE6uGV2DccPaQeds7a+P/m0
WJ9kqMIGimZJO/lSS3ezvk1Vh4pN5sQASGHi1zaRQuY66pS+XCwS/X4bexXukNwB0tK91FSqJouv
Yc1WMgmIPQx9jC89N53eVQUHdTX8JbSR1jayW1jWWTUi4Lc2v8U8Wb+DOAgjfd4zT3dhlBEuhXav
D4LiK9EeDTpUhhN9Dg9HwbiPu0B8Ou8S4IK3dcXCId/hG03LruJFZQN0gqJ/3G0tvE6dbEfGaDfQ
JBu3U9CcaF4ECynAIJZL2sBeD3O4DNm8JrrA4v184w91GceFwRpyjSVJHYYherK7fFkrsZAtWy4E
55KEueAY6purUmXdfU3yevGeEAwbG3UfRYRFNUggObCf0ghPL+8bEd+erZr3/5wbQC8ogYez14Rx
qHuHm9bMEP/dA8umfuywjJIR+uYBIyoUCnbnZDEiQZcBfaT4Fd10IQlSGbQtyDngS1Z2T/24OFI5
mTNxBhNEgK/V+KStskGV0QEE+JAPVpYH2dDcf6RVdfwhvw4HKSZf781QhMDpAiqVKhvnEpsP6Hox
A0DkgFpNUwr4VBmxzzaGMt8CKPRepvTR4uLvzpyYRmqmjsRVgqVyvOCKmk5daSRWE7jc8TeOywc+
S1KNZLLTzgnYAwhRcl7oLLyx+9TwU7uZJFSOscj45jAk0hCMM862Qdin4/IWxbDt4j2EJpsphDGO
gAxN72Nz8uI3gaKPE30t0dJhBTlMbV2SdzUKN6kLyFSn8gr4dZntkFw4T6lQYmGY4hsrzyKSA1gV
RcFlkeU4BXxFQEd7p64C1ckEw8LHrCiSQFtYdk7UlyhgOZLZ/UsGGOmt8Y6Z8vlnOf1fboU/oG5f
L3fh0Lqe1mTcKXcsZc95CfABavmQhtw0x8edu5dxIh2jnISxwlJ9c1BxXttQtojZ7x9l7SEDYGn4
pvzCjTKmdef1R2lgH3ttfST9D/8H799gT/oqR020/G1w2TjB9De1fzgj/OgeD2U+zdbUgWgVSDRw
rtNAEJKPlFggG2+QCv2lcvekb0FNyRXcAJRDVCiP559ddZgZ5AB4AYAJRClGtzKyVYTq/ewrWoKF
vI/Kuwk9i6eacn8cBPAl8LRG2Tm6GIld56CWHEWgBypZdKqAxVX0dqPmRjAqhNmS3VoPAp5Fe5Cf
MWZUAUTbxbh2iCrvY6YbnKjnTq8z+meTYvKNY7uLmN+zWB67Lxfm19XlTOZVHawo49AGBiuEtgp5
GsPu7Ggsq1Bq98cgLrpEO6YgbYhivt9U3f+khhFA8sYzu0X7m2Fwv8QDj50lXgJTrOg4MD0bxmD8
CvJahuhLaoOk9AVEdAuLw8kxfpUbKftGFsrU3ZImGsTpBo0xKCpCzcmV/WQLnmnCGKFgYNtMQ0xq
2DPN/0ijL6etqQzxabbSpWM6IQDkPRlz1IdssxxGKn726kP743QcoypPLL34PKZMrI8MYMsDRFzn
7uF3XM71Jl924s4B5LfivMYtPZP4mc4AxkYY0RxiARqhgYdaFPI97wcmt6NBmkNGP3j1tUqjpTbV
cHLvSzUMZmvJxssRXeDgGJAz4BtMY/n9grPZtP451x2vwzF6y1wUbpWOJF6hUNhOhlkFFfl7Olb7
rpJYUZJ2Nujd7RbmMN9CcAJgab4cDw5JjmvjZgODCFfzkmcojBPbfHb0gXKBIa8+uU4jDTCuHa8J
wkfzUkzk4Uqwc8gtH5mDxJHETmpJjPn6kKfeZjy00R76z1h3P5WeYwKcMWE1q+JISIMetdkYITHo
e7dDLTsPEbfBmI0payNR2wqiuHD5d+Gy1r+DJg7GUooT3xlreNQU9B1Wt/WNVbZIHmtWsU+Z05Qi
p5Gwa290UOCHceY40Arg2m0ctLhzQqvSLjDzAvjQiuxYZ8ydUR2PnBuSyBWziiap9DU72kH/9CIg
BxtkLAQrDuSxExdwI+1dd6FBZmE1pvLdgLYdi/PTO2m19F1a8xn3IeURFVGeL5vUl0vsbS91ZZQ/
OpGHqy1C1WrVElfS/vu3LqAwZuZe3pY3jyPSNh2ixGgFc2FPLFD5wEVF/Riq1exKpP7CXv2rdOBN
p2tngCRVcMN1MrN5v7JEo3w8+SKenGGch8ZK6FdfVLZS2NCBUQn88q9KG/6l/HtasWcdJyL+HtiP
w6s2711Tju7Bu7BUcbhYa5PyyW4ooVFAMdNouWRO4uftFEXU65rOMBfRfkGNaCRzZKp4biVhjgmq
rA00VAWXuUkSgd+a41Elm7eg5tpvO4Lv1uPf+ZVLG08bGR5hIVsk7goEprun4jjvsQP3Oc7E5Lyz
4nxV9N0LkxWCmH58Uv/LFJE151MEskwOOi/GeGSn2QAn/7k7Q+EX4hoClbbu1S+zNISrfu0sYdat
jCmCA4b5V3YvjymENOb/XxZLz7pkfumzr1CLKc0CHcAa3/KmiMkx8LpCp86rmNFgcQuMAZtQyjY7
b4LKx76le/DRmGDOukohWcGky6w7ptlA9DDqycEoa1BS7iT8/ZY0uRnsHrNGsPTwcs8AHkxOrHue
i2EWVt/hBdieTAgaOMtbCKhgqGrwNIXz9ffpvoQtkHLqEMoJYXbuI7w+eu3ooeWtuiTTQaEaxAei
4W252yzKzPfi1SvcVNH1z72HBQgN4/nJ6M75W9KtKztQoTAGH5zve0u1lkg+a+sKZOCloRppAOkL
yCSeRP1BA3yUvdqwUnpsuM4ruVlmOFZX0VOJ4Q3xM/K2Y4Jr8jgHV4qrX/GpvbiqyTdH5pH7h+WG
kVxmuliCPr4HVIZPffjwaxE620E4XvuWoPn+qVq0Hn+n58ubHchh84UthLFzvjuyA638H6Ud60J4
R5okYg/Hsw7WGSkLtYKbo1eO8HruEGsfKnTkG6/zjk8o9cN6Mu25U8Bl0T54d6wJEq9UZ2V7WuNo
LgQD31pLXyThJnWQ/vCRhf+nV1fxLQlu8NKCb3E0XBdtu/oHGK9q9NtsqD7GGNylmNBEMlW+/eV6
6BGoMUJbpySwtrs1hlg1wcZAfopKSHW7pIJVuN/3RmgOHN71YvVO0zDmwRq9DrE2iK5L0GNgkL17
cwnABC3SRoc/nGGC5UbZ8dtgeTXG8S0wUKO/dXwIkOBvbpYuKzAsr4xqdRLCpWHK0S/RuJPJG0Ss
smfv4VUyH3PodnT5cLekEWj8oiW5vErMo/jsw/SaU6oqKXaMiLwBaUwGND+olRO85Qb+TglID8bm
u0X1UX6FTJ8+YG4z5YxSKZuCfeM18UgJ7uLvUnEzPCJy+klf82fv7BqRQ/lt1fxaettI4QzRdfJD
Cp1fCq0He5P4Cz0ig9Y5eLuXNmLTg9HiDIVkTG7OQqCbRUyU89ZoO6UrcA7zNyRPRdpuMXk3Par8
Cewo86a56gBBm7BQX8nfEP6IvZOQWfMqJTrQH9ICIGjf8RJgdttlBwpwh/WWdBB7UN1IWLuEwjM3
rWA9Se5kYH4bXTtcLLgD6zPskVc1HTqofFZ6JEVQMX2mcE5mlF3GAJi5Qxg5eCb1CTmXstHsdqVa
mSaqzZugJgDtYJutH6z6OmfUyY6LObYTc6ZiSOKcluVMRCnkG+MLyefh4u2oR8725CgOSKx0a7Wr
J64KXk1nnmnHafmNIzBqaEJsPr+KpzzrTJ85+q67rq1CL//nfOsAQ9luNTOv45UJs1bfO97PEomc
DLzg3ASkdjUl0rgwiBn8dL7AwdQ8P0BU/SRPFOU5CS28j8GwnP2322OXSu3CqGl2CqP53z/nhHtB
f7inTOZgdM8mfTN4xCVYxVCqa+hyZQXX8eSBZYI/Rzzebv5HBk7jBAOkunjIbTzoOI9+9oF5bEux
/lH4YroKXsmAVZFd9zu1X6g3iToXBsN15QswbrwyMkE5TDi6ackGmjwQkLt5vA4xSGR/DQckNO0k
DhN/XkQMoe8twrfsEnGnUJKadIOYkT2irmDkyfCmwSduaFr/H7hIa7v42QGNNzG8/dSV4FNrNLfb
Ea3WBXvItRrgi08oIeeWlMDGwJZytviZvgv+/z2EqpQNcO28sjZbqyTxnBqfSXmrUNjyi+y1r6oV
Nd3Q5st1Mrs3GSvfx8sIUGaA9ZLNIh/XALKITezYkCy+QFqThQ6OmJuhXiHOMI1xKQw1wiAT5HAG
5f5bGDFyQtlyYdOijzsJYs/cG+XIgpw9Tk+PxDvgSqJnyWYHuC6oi01GsPRDP+D3GaNvBjPKGtlu
01oRfKkTowotKSvjjgHyPRcXDWAX3uJB1goSEew5LKOT7CNon9a1BdOG1i5FC3jV3H9MS9crmi9W
VvvIMLACxgLzN8FlqxJxgPD5fVhz5ydrr6X/KRBKE8rbm2ZpNJSI2qPFiqmogiIfsq+O2C6uMqVf
yVpe0e1eFKWyMLDgD9UuqsYk+cEby85nNfm0GjXW45BeB1qgMa1BYy4PS6Ur3IkzIV5n3Nj5OfAY
EXMnaFqUXTBqSOq9wDUYbtIkO9ShYNwFc1zQYdqQEsZW873LG8hMMBdVPos7hc1wDUh63R+8SZHs
Zr+c2VWv4Fs0Le2SM0wgrj5cWosc1IQQS72PDrq9JCH7uCeCeSBq2c9NDrbKoPdhLaSV+A/+Ks3V
ioLDJjSht9e1EG5y4WDEPu8hquJFuhyKQiSEEjvJGfTyO5qI4FXDwv4xbjPzpDJ00SfFTc6SHmsR
aM5UZDMUTcSoCLQIPPhbKk+ja9U+kkU7O0Cr7BMDqRIlUBc5uSquVVkY9Ieis8ipHpbff5ibIxtS
TBIFS7Kc/UeVFpwlLHVpMZxH5uIud8vJdAs3jBI2hcsm/ZplBLcD+hWFnENnYgAMeSm6O7i1WbB7
CdE6dURBh/G9yL89FqJ2qfB6UtXLFsLBHA+kEvsZrFpIsim3yP9HKcGiZ9SvaQmAkhFkdRUe8Djx
WhxsEhRyqFEqpyVJIBRfeB2Mxd36R04M4vnsX57Y9yYdWLbZdydn0+TxrwqlF9DpX9rDKxap2O7a
U0kgDXHl2w4cAnRu9J6gdm20BEANEC28HBeWc9x9SEuBWssHUMNAO3NI1UeHTTdSg17SC8k/77E1
jyHCwdXXzzVik6aeCqKz10t8w2WaxtQFG9Y9oNSGZIg7UzR6nRV9IMYISjotHB7m4NG9dr24AeSI
oWlC1cBaQd6JWneDgT9A6vXata7XqtHc6f6S/LioO0C6kDUNd3Ux54QUBE0i7runZSBjkwqljIBr
IDfWAcolnxrCrLDjofvXuVj9qS6mB50CDLhCXhsB03i/m9x4rSOQdfdHrxSm7uciH84tmEwqzxfl
djgQDcGGJTlylX+Rxlg0sWRuJ/XpM2tWkIRvJ2skqWVRHAee/cK7W6h/51j3bpBGBXedNw5+gFum
JzfcG1R4nQzxwNBpw8fsJM27kszJnmQtNiULopjhvse+2qe1X/9CLqdZ55sj/EGIl8LRfRBiQfBM
29bYskQju/wwrCD5WplTVvHkQnBlnFqwBS0TEV85TnaiSTkOD4sjDbLdKzaF3H8ArX1rbBftBoDX
8ix/63BzMzhcUn0HLK3rsd/ybjTYyVPN1yXLfXDXIDBGsUFuBHoWrZnmwLE89i24cXfBQnms/sWg
fSm7fT5wyJZEM3H3TJyURW0GnWCiWanqk7e06HHl8wBZg61vSUH0vynezRw75VzVm7LoJWaonMRZ
tI9t3bYMCAAVlXuBZdSrPzmSxjRXN3vzq9C+DofsXYwnzm0nz1hn2yyPFgEJpMrybR85S1xUpacE
J5JMZ5cb7EL7bqjdWJRph4czD+7W4aGUg2/PoLoEZWoyJ7bh6tMpTB5L+WAxyJkj3bmr7C22pE+g
KJOV+6znKNg7cgkIsUWCFGm8vqJf1ArdTgtGU2uzCgP/paOAxtBV0bZdwtTMhYH0rC1/I+z6dsem
c2tuBriSGRRqSBaWrDZK+/x+hscLhUigc6AgVKduelmF55m31uSfm5EO0Q1lkIIwWLF66QIka/im
hHtNLCQab/O/HaVOeFlZ6i19958C8L2H+wT5oUodRrAlJ0u4/8VtzfbEneZowWGNAOgY19M/KHV4
j81MTIruymjjK+a+2sLHVxqSuQbRVhUISOWdMoo4fMhh7QMphgFFHcTwd/KEW6peS9pkWwaFhSOO
xlOrjqj3xUQAzKmK8sH/BL7ST7n3C2i5WfThtZRlubolOFd+pk3weXmQ4oAWm0Sz1z60a+qiSgrc
s0J+8NGxb2ctAqZg3mPPFgfP8Xp9qT+M75UNLZnn8IgUvm1YE2O3NyaFGPrPxEwnz9HjV6k3oNg0
d4Qqgn1gCRoarLhRwzhqk7bVOqTRTAYH06qfcEP94/xxJ/Hxz0RynrNN49Ut8WkQOe3xkiyurG3R
DzjLVBLlkOHhB0owrMDQlo6yN1y2w/0upSR877wcJPrey7/EwUMx2EjRJR24jtUnBil2m/vNrgks
W0U0HdPPbpDY5fPZpziu4AcSfAFoiWz4x3cNwa7pdOhPxkER/u/aH6TPSnelTEEPYoq8aqOuIMNv
reYCOJ01XwU2IyYFzfTBMS6PreQm+dJqY/OEKoH849LM6WGrEQj+pnK27CyHjAObAaeJTqUWQ+v2
gD5ZmFOBeiLZ7j20q2yC4/1Y0VjxX1WQ+24fHqvKRFIjA28k0vnghTxZKqiWFhlIT1Oew+PGih7+
wdrLn97+3gNpvgZGfDrQhAMOvJBGv9gyy8OldwEOHIEU1VP9QuaHoI0KcMJz+d2mR7b2sV/MJo6A
aL8x2yPsTgM3PEB58Ioj524C8CH+0KONBggPSFsyaXisNE+XeD6UZWseTgbO0sUW8aetQwj/mpRi
VdPimlmqGUS84vQuWT3q8iqkHSuKIv3VC3QhnPQifda46O4eupDGo1Ha78f4DOz4kbf8c6V7FR6b
jdnEzF/S0etL8BLmMnEnersBd7bPEO1YrRVqWBkIj3ZGhHziWvqjyNcmKCMQ8YecPh+DmNMYnzJW
VYcNIPn0lk0K/8ec7CDoO5iG/h97CSw8f50X9Lxj6s7zsXlEdrcJm2pLzw0MOEdUQMIh4/PXjPcP
nQ66xYcrEDlDCexOqNh83TTB8p47z6Wr3Dy48x67M0MiQhv52AkCOGjku2IQ+KP89ed9yy1sko0v
77tyWVT5622VtwA4zY5X01j4UC0v609DfoS2Svst6hFUXTF+0wZz1G0hCL0NSKrsVRYWCHnXgUnX
ucGgVFc2kiXghV2/wBcwy4VNJA/zxYSIN1KW7nKgeycLVR4S67yRi6u/WzMsNQZ/YwprZl38Uh9t
eDi84RwUTNspfly/obv4DaDEBdILazOuqd2G1MVN7BEfUeKi+zdyMAlo2UCnq1iU0eZsQ1YipNfl
p/vCtjJYuik2/d/qWVSITPRL/U9nrQX7MkDCfYZ9ekDjBgyNG3YQ87BypNdhSnPhXr6RfN1hD6Kb
QnC9HWnU0sNnA3hSnwNlR5QJbyiA35qO/Qy8SuKoKQsxfyi43Cx+A13qH9iZ96IZTrQB4HgnTY6L
ktRXIvCh9QFkAOuCmE26n8/x93/5ZzzDGZ8JJgWf3u7D3EliL8gi4pqyonnPLa+XnBkBHqByxxDJ
3f0hw0oB1Q3lkM28kwKt2TN1bjw6f6dOCWjnqoLd30LHd1MXmMhFF9+eUM4SnvQE3W/PzOOX1zYo
2kbr1gBRYCsb72Wnqs8gY18a9GlXKcixSKlrexw34ZSO0B/ggNmxBmkWjEoMZxZYXvQcdC/yoJ8K
44trRE68BcAV00boka1V2C/8C8JnmmdluoQDQrokmY22/cvIDuPsWSyeFiswJ785OMQ9qxoiZFt1
3qbkm8dOfRcQ3G9MLIdpVDJGSnN8430G1S71hYsLhY3spshMf1V19ke95xhymiN3O27hqUMKhxuV
9nEH7VugvELLaIpaE3QjGoL1zmQl1k3+cB4sZpsEid0MOJlZCn3mRuWVPuZuwjDP1YJ+8PzRRM5q
IZVUk1lFzHPmFySievUIv8giA8pEg+DU92jgcYFAhJPDwfiyo7NAod98NUq9m939N23ScRUZELd2
S4lkksYKfb8BaOaT9hSX1yjd87gf/839bMFEudkyXZu83f10Icp9cn6R6UjEz2+A024bWpi4EIOQ
SRc96mtIf2bnJoTPj97bhCyNe//D5y0PYcrus28o1SaF/bWCdA0ROR9EnJNtC7Fsix7tSb7/jFX6
5LQUP7chEyHKhjUm6Xzgk76ypvGU5cjVCGG0yQFdSXfYchQXUJ/wcX65wkBIwHuoluTJP7peerOx
HMPFfD/W9pHGALzc0eV7pJIgsl7/k9HCWlRGPxd2HBon4cO88z9DCPzfXrHj5X6MzXZnQqLHphiX
eslegGLHIUbq6VyrktPNhCdZa+/WFydp2gza3pscw3ToLKID87kEeaMPICJFJhlNYXJjw1P5QOXN
8hDSPd4KK3uydDW5lP0RzlxCHjZwutLoa/QYXJW0cAXLcag1jjR3HMS6TFNqeWhpPedW50fiZh2o
TGEEiO7i/TAE/F7ilIO2fsFKZOBfa/8UrSkp5g1fZFoxhBtwsF2h31Ousv/2LomieCGXtgzv6pW3
1kh19d9WEi+vcREfb80ta/iowMnWX/9fiU4VzPCbv2EbyJ0JvNoEHBJzDajtp2UVZv5Ry4lhlGeV
QsgP0j4S63Ucpw+hQW2ZufbgNnWPbLPHDW8g+KdparUU/A3526TPiyVyt4mxn/fQ6CQooNb+ON+Q
/HuXGyh4Sg3QwHETMoV4lcqsg3RCnkree32yEQpYxiBBtNjsZA8hzAeMKtLfQN0kDHzG4+wPQZl1
IPE5zA1yV8O5d/XOWT8GrRPaSyDJZRG96hhoD4juAfcL5u367+t4bsvE3gFDyJa2NG8up9mvMzd+
PecvPrhY+qYAqsgY4r4pscyaJyr/ZShSYI+fBLoE8HMmeb2JZOkePEtBvLd7YP/WvFDNngy5m/Ha
WMziWKC53ZXg7ccsRM6HMcwsm0iZGllAtDZrnZL2J7n60cJy6rT2eY4wiq9qhvavKkk+P7eac13F
PIKh/AzaHPcsNH65yZ2V0c08VnLU2PTAvR11GP/zD0R/RpM/5qDVtsKyxgld+7NCIV69zBViFsgC
bsHZGTRNgw6NPFUJyK0/gyt6WkNDcYrVvsLowPfiZnQvdUWl27LJdsLyYka48O6hlSxdcIxfCirV
0+Bhm9PswqSs471KlQsai/K9yvInQq9d4HSNxS29x5uZFli/7OV5BVA5r1+20nTAMTK6K2y7GJuG
3Mv5uU4m9YX+pROyn7Ea6gFtQxjml0hLpspgD5HbHBawMAvp/qQNwZRilc3s/POn6I5NlF2wb7/E
r76Pi/fApkC3CnpOXrUqgEHxQN1FqOBCEv/E4T1Xc4rhh2l6yUIlZ5cr4bLmPLS9wNSKeBxkEqIf
KGzTWyZiHBgRNKC+nKkvb5vrT+pQghysRCTk8rFxwDO7C9Opkb7JPexVKzcqm2ENXhPtkndFJA/3
zVMuQ1c/UYzAzWWywnbjxdDH5rWkPHoC5u3BsVlmUSoBvgwNiyfAzE+oS6U2CCWOzmysVISPmf1e
+N94NriQrQfPBc5wye15Oa/Ez1ISx51O2xKIscgmIbaXeZkQj10hZ9RS6WqN/ZnFjRHW4mC8Vqzr
CyFnhLZHojPsFwZ3ltAKRA2Nl/kTp2fy0qdeM24cKFT4YgCP+B6nRF9GW0GQctNaxKir75TJyk4L
0xMyaKhgNqXYEPVot5l7/tLzoQS+L+9YK9RGx2ODJaUtjUg8lc8+faNvXJyKYMmS4xW9KtFwxfTj
Y5MaU2Jk3Cz4o4dj3AW0NeIpPMBnb0ouJarPVAYGpzUsfLYGRGc075uaLqlAgpsf9CGxSyjfsZvd
kziCtdlwrbWnYn4SvZamTnWJafjHedUQx12CLdLEPKee5pj2VoZ6+tX7cWVl/LdheO6DnECGM3Gh
muSEJ/hGySfNV+i5wqT6bx2k5HOnfE6TZeVtbABY4N93bZ7cPgfSvYoksRoZOO5awx88bjTMmgY2
tMmxJWe9Fsn6/BzrOmvEIa6NXFqo3u8MUBwUIxvywumFoq5ZZ8DNM3jfkecUyF3IJGkO/5kn1lju
2wNG24pW5GzMDJ1ftGP4UmnbiecgKH6V1+F+V2InALeEmupAP+Ev84U5zYQcETlqz5aCL7pgq+0h
XnMXnXpQ1SqXCp4OJ64EdxxZfDtqK2YuHo3G09pu+temhOk8gZkN/2YF7zO8xZSmoaNV0LUGwWEP
zJ5QoW3nEI/iYrKoZE8bs+cVweL0PGq9zVTK83x/fNpdjh3+lAtz1OdfQ9+wJN5hTtbz3ag6n3Ia
Qx7VQCYP6sG0JgIJFepM9lQsZj/gA/e+bIUfe+tDfE+QsWUHecRXn4z3pYsq8OkSkdyXE2dgZnVt
RGzrAcvNvXp30bfA+IyGm2Ft/SRIu5tqxcVMpgG/CiCyIPAdRUOgIIMaHtD2bQ6R/h9heqxMYRo5
uLuNDh7NfWPilJ54O1O8fZUnzZbMusefpi+qB0gB7td5SQTh0Wg3nHgsS5hivLjxfY0HPpaj8fBa
7RHMm0KVmiYxjvWmaaNeqGAvw1LKB/TDSFmt+wEMdco67Z9sh9Qej1XMJTuAt8BND4hfW/CtrdBi
VUDptGQa4Jb4WuyO+0vmillYuPuhBxG4e4B4Xz2g0yolcsFMkcRU0nbi3eALfH/z1dEIEFsdzHp1
MT6vFFf7vWYARw/T+F5sJbA4XMgS5ZehWjuOVLD/Y5WSmX8+EQX4/bNQ8DUl6cWoVBDEiUDNs5E4
xYNOzeadmHxfPSyTG+ZWhopkZsek/JKhHbSvMeSYZHnLLE3bSxBssY+mH4GR8S8iaLVU0X2ASrNM
gp9Vwi5f8BMqpzRI3rCNOiSvpWHj60Ssh+PPrPs5Z2LSTQ5FFqnsdCLWUGH8zKB544HnRobd+dAH
WH+mXz25KT1qM3vAwf0/w+wITt0l+Go9Bd3xM33vG1A9Bb7pd6OyhDuQ8VY6w1m+zFgV91rd/xU/
7QrLIPR9VBgoy8TndA3TYuWo+AYXcT8xMM4N1Bxri0hVNgzHLx0kjp9jw7tY1xacp1VWS821UAV7
kLvcA/wOMXif52IfyIX+1IBsOkwfJGpNtH1ufhN25sZsj79O5WiouqCDPwFca8XJPcs/Ks2d11FT
60VeQC/IRC6SwrKwzlwSMQQ1KER1EZigQc9kMoavJjhLKPBC0v88ItVNoIBm0QxGu2OxlbFcynp6
ZKMPr+5cLpQSc+uDExGvAZPLeOpK+9/udRRXEJNRhKAQU5gIEPNbP1Ap9rvrOOeeXvQMz4lx4RCh
hhXaayD03oOISDWOIeCrT9A/RAdCeL9jKZB60Oe/3DZCRBU96Idui++jGQxWmUELMqS/A0+Wl29E
R4xqX80cSzAXuMRqXcEvOaragnk91YwuuHV5bOP7r0HVa96hoShaYLCBLhi9ZWDQTAGuSsr1no9A
m90SANE1xoPqHg216XUeT19r4pC8uEQG7duTIaR/IzXjQ4xni8YTpC28gPEa2i2lv/IbRY66BB3W
n240HGFfqLMAM5g/eE1bG0QtozA9kfYIMjtv2f0rWzXXx76WJ+uxINOm+aG8N5k/LSkszH4MdS4r
hhTFSAc/v24Clk9mpl2krFbXM91P3cagaI7dLMzhdU1R0CkKGO7ebI49k52ORbdUIjeNH2DpxDBe
7prXDMt6vc+H4yG6Mt0YZp0OsmwEcM2qjyHIL3KRy1hVB4bcTAfGJF7e1yMzJNnlE8ZWVe+n9rKD
hM3+Z24dS/q2CU3oc2XUKHxtcvcblj3m9VZmcHdQ+096KbP8WSDDz+oliGBZmXVHqdIfYKf7gNVI
3JhKEXKJIkiOpDRuFOmlaOsFIt59FrroR8k2EXvoWODVJA0jAdI+Zm1/YJtnV9O0VeZiFRHExFmK
2Z9Cmbomoumd1MzlbF99YCUMdTpxeF+7Hif0nsnaUVx6xjHPadYoWCte3vIdZkKJbuFIPeJxgY9f
9yfYRhewbiJS9VvMEoE4xXEH3nTqJy5Cb5plv29AuAIqQIEyYRwuNDESQAeNURTMiDyRUiGMwchD
dOnArzdyWR1SkV7MEKuLOkOwjzCjLSm9hifFN/9jzzXxrXLsGG6KIte0lxl8iR/Lr4rSSC4Wn0+A
KMh5kpvEdftsk3556/azPeGHGMepcggMSA6RD+WjxVj1NAcYjc8F8zYPwFMgAaKQD3y5hWBpX3MS
g4g7S0M0dKjoQ1Ypy8mpNrN3Lx6I7vLaU2SdtXTI6fXrcspKp5v6so+J8dVhc7Rc3+A3uU83icoF
0SGNRyoIhlR05i1jEeOT9d6R8/ow33//a3Vybx7RM00drG/YViVin7IXCoO1PsLLZ2L79USNjsyZ
lNkqulMeFXLT/po1i63YSg5M4MtSReya2qCCluhci35uChH3czsbwNB5itjrz3rXGBkpNrM67WJg
vHG5hoYTE4w9cJKuW8mkAElzR2JRW69hPZNIFOzN0DF7Ma47DbPtkTaDenUdusNfUEx88HfjklV9
DpIoKxLaUowJI7prLjq8ntbrzst86qdfg9G8jm8qemOV2/GdIwNwSkjqYXcXjnid3dNEJeVQvts7
XyEMlApEo1YJm2/hEaq5ZZS5JEoq+xJPjmQiDUTwHklR7tI1ccJ89YnXitO3uKEc5DDtxVJcukZN
8Rh791EDBge96nVM/M1Pix3Y6Ka6YzNssVQGa5nXIMChCqDBSNSK6aMEJ6xV6cB6I4kZ0dY2tuTs
Evl5lgI7sTM10KAVL5b4kwk4fPfM/tYKx1Pe4L8pbW1bBrLH2PHgUL0Qw6EDQx6YsIeBEZb+tiYW
vlqD6QtlJDch92JsOFuJRCOU2ncn8F8/SiLleYhDCpPik09Qy7ehR5wxmAa6vrPftral6sRRM4Hb
/Xlg9azmrRBy71+zN1XIu4A3k3nK4EPOUpHfqviCJdQwzvi80TKX0jf5CApN8wywknAtM9HbLmw6
Y4RenQPsN7d19FJ4neZ+lcCmktwoKArYrXpZ1sNAL2bkN83VASdzUgI7oMfchb52STTwaUE+qhHE
cbhBIsg0wNmJecetc48ODxig/qyO1DKPCMzM4JoS1C/KOJdqsFHAJah2wIcj8fCMR0MLx3H9C2yJ
Fk2N5SnAjUGUjyn7luGwpva54Zr1NdOnIj5VUkdYDyvXd5QbMx5Ds/Q+QSzPXq46FuAjZbsu+3i9
K4gzS10TjuPmSIzpPPXXUBYf+BcYDsdeANEytDHnQe4E9LcZQxTinFd0Qb0t3vq8zl/31gbUnOGA
+g5cLXtzVKXwH+TRumms5xe/7ae6oM/ocKDRAwV4Tq8UFI72406DZgsySfHUpf24Gd9cxeqdE2KK
FYY+DQ+R3wjXIhd0BYF/ISH0rOVQm4MwRwKBETSCx0bOAf/OyiHylC8RCJbExoolFCguUaWsj/1V
G983MKTIWhoXFlSXoMFR7V8U5duBelEqLYeM91SQGYWQ4BqnY6/aynmK+ihO58SFKHZB0CoG9lyW
lgMlS82EjTUSEZcIXqjj5jZa8hj0agMAuY8yugCjdCCUxAnV9RrtWKrZjX2R3i05HpuyS5Y/0OnS
iwnZgD9wOMwcAPi3VXUZPyR687bJrl7u6h0sJhHmiCW+8/lSeCDR1wEoWCpmxiSo/MUghb+ap0xS
uPJ+z5Tw/2BomnNpTEbChp5CWBN+EAzIAmclGCmWUOskVhNh0EnimAHWuNCzbNGG5Fx5yEiixguN
Jk7i6m9SBPC3yR4Hv4Uxiz0J9/HYTzPGuP6ddTdhLESw2UmTr8rmWsp3d8kxBmDNTvlyBAsIRs2F
9lPHutwD5nR+cwIwEh3Y2vLtpjSF8kwcyfUtssXYUNadJpGPngRvfmTsWBfaJcRol3tKW/L8UzN8
0pLIOYhQ70l6cD0P+dqcrNlRJIuR8D8h1nLr1QTY++6JY4rvIlgkbHWu6r7Kv68nOYInkS/rY1U1
IDnR9vOIP0XxQIEdraYvBx9BUiLyj+tMwhMBwcuR//aFH0B6vPsmlsFj5pASLA3MKxyDnLcWnv6r
zwWJ6afEQZwafcHTYCiKT9PyC/Kf43DbEKEJdLGiZ/px14dGFQoAzx2wto7TRsRv+QNDFpFmm2xL
a9wucQdjD81wbDbNqkIrvQoyB2wersoM/O5TMClu0JCggTwhTjooFAQzapYkkVU7zS+FnCM4HplI
ko0WGWm+cQJUaNOKZFUbB7BqjMp+1pOpJ1pZKvUY6sdgIRtoOdydVvncWQdE2N9XYk9A0JlyHSR+
1a5N38WmLR8a+Ww0iE98Xhz49dEkurakcEsj5ETsgXtquXu+GM0AhpA7pRRip6RtriT8PlsyOU1p
HwOZCmgHlK3fGl5CFEPcp6zlhuTuVgqFQm944GiPewBBLMJHtmiDptubrd9Rjnv4IJDO/jdgK5lm
ivZT99kpjvutjhuYCaIjG5VX1Niw7OPBqp2H9s9jrl2TZbd1SLY+tSMHol3ZNA+whTfrriGp04lH
sjB2rio7QXpCQzSC/PXGAhN9JG40EmqWmRNcWI4faO5DPYhKuNWqz0boMTBoXbOgvisDictgWPcP
V1t38fThjYGjS7ukQE+pMllGH5niZX5du6PXkqhR1N4uj51wq7eZBCh+oZqyhMH3bQSMZVlO8ZtZ
MYEYv4jGxTbexeLwIB+KvtyZLHaXhCpoZtCXOVZMds095k2ha0+9d+8QUDoKB+uCwrsyk7pXTPVV
OrUDFVJDjnMs3CYBVUorY0RHy/lCDDmItzo2594TngD3fkJZ+QgtnDJQH7HNq+DOWTdFij41Co82
3vPuU2UiaXqVC4POLPbmQ7eem4a5Kb7B3XBgxxj4m/dpwFXCYtsDV/rqS5TOJS9IammoFS0KUcnM
r0RiH2vxbZFkJqTWeMpE3rP81qpFGSzJoWahEr1Q4ZDkF7aB3QQPuKe+fyoCAviv8sQ4CPVYy3Yr
0egndYVEzVlyP3zeruUcbYJjegMWxSe+rgiPGdC1yf6THXsKpi/TIaa3ZtfLDvNxT5jg7ZTDIUvB
A2bU7czZI+hR6SF6Yx3ANVYk8BPg9zOtyunSHUVjC1X/1OOwAYmYxJ558VcT5UDT1SzxTBIYHeVo
2+uowY9IToBAijp5iuGUBt/u0Rg1GrwPzBNqku55vH7vAt1OO10AIHZSCqSF506JlaHLqJ6r1lW4
MdYFsghkesYT5IquKUwJAPmihU0gip5RXeJ1Gzus2I38AmHdt54dR+xRtO3I8UhIkTpwesNpTAQ6
44daQ4Sj8fxyn7yL/a6767jp/E/sALw4z7J9ndqpf4qlQJyt9qJH0oCF81Vd4qem52pIlJ4li1rW
wS0HgJ9HGe/zKXIqy/YOa77vkN/QV18Ox6+x2bNjPyZYaJQL43vPOFpjHjb4PuWlRD8pWvi34MWf
ynXeDa1AVCCPD3VsP137OodcSxyzqXGl6P0kLy8OGPPje/IP9o2hoXsDm3VX3vmOrkdCGuU5qOVt
C9l3SQluLT4Q2NwhBdTka8Af50yXVf1b/+0PYpTDi/cQMMw0NuZR2QW4BUzw0Ro+gb8RSWZzZg6L
l8VFbne3IT6nzkDXGrq53C9b+p6YKFOtk7+CQQMGBkrupGaeOnNrAhGU6TfLHkda5DNdo2KseOVW
QY08ueLkQ8U+d/0mhFW4jCpcDnI1BdTP2yK3VESnzx9V9PkxNl80f3S7bzhAJXwJJzrvfIduCG7+
8GMi4Ahzmoaez5N0Vl2Qs5WQZpaV11BXts982gqc5sTenYWVYiRpIJj+hIWprjEmvJD92lgq2Id+
W1Y6XzNo+2O7diJ5PEVSIUll6R7Y/OCrP7zBYc3PAiL6I8zVfM+Nm2fSNx1uTSafn7XpCnD9dJzu
ELeha//fXGXlQnFLPe5PUr2xvcmY7zHREBH5+qfH1YQ94LMKOkAKjlzXUCbf3D2mdvlSdUs9nlAJ
eFaF4284kGZFubG43YvJiJJ5oogHihFOx7B9gwnPat75N6TG37NyC9LFCaWc6Ku7suShmkktDZ/v
K/uV7bRnGEeDfglhGsrtoeGvrEeYXKgCX2t4b9HLfQWc45TFlAzNW2c9o9FWXfSlZKCqf+BJBUEh
WdW7h+aWj/Oxkx9Lpd+5ODZiJ+1h/LtPz0U/ZyQzRlkv+TVUpFUt4uetgu067qtUYjaIdpt3TFQ1
jmpEotFvpQ0UOvceNvWtjjeODbWcXDPtUeZ2ooFZWcwPn3IDWAC04WJ0HTrlj5IiVY25Co3Slj3C
2P0sh1Z9OBP704m+6NbsmmZP9tROXWDpsRoNAAzqvl1Kx24XhOO7yzE0Bjg74DcMZ8qG3RVNVuzY
nP9cAtufrgJoIHXYsgKSMjiKSvxUi2poXt1iziFtfzPw6B6V6Q+K0ITUrb6QqkKp9hdpbj+/rC+C
mCJClPaInK5j5PcsFfUv8JLDJVvQ6hJ+5EpV5qVJfZR3Y/tozzU1SK59ymW+pLsQEOy4JV5xmufp
N4+E4WFsWULcyoQUlqwMLZ5EDwvzvgux7BCekCIVxh5WVR8XgRrhoV64nGBHPVWI0XjSf2NTu4jG
me9wcnGtnBUmfTOsweSpeCm+/wlKF6OG7wR6uKuzpLq46/eLFzEW9M2lexJBvicexUlNoNjq/4ID
1qCQiKNlcjR3Nih7HGjfH2bFuDzPGHn5t39XfRZlXHt9zQvtAVq3rRdBMN75Al0zshYZFsanoemh
a4mmy1IKc0WBoEkwTxTYpNcpyQx+trk7Lc7MtF/Dih6RVX4O+T1R5CwownAUilYDMNgLcuS4IkOB
njRtjwQE6kgOZoGRr4RhOOFM0oZ3Ja4ftzUhflJ6nUMcq3kXec+DmCyh3kQLNWCoIWDBtUUI18Ah
WYi0F4g0tgxOnj8NCC752JnsTHPZbgY5SjHovtQvEO7K5hG3CvnLj09wa0w9JeHQ7pqN/vYvSNUe
9HzSPm0T1bimk4Nzq3iopFp2ZF2suSF4CDSmMS1EJQ6ef3Hw2hWbLP9qGptUGnico1WOHd+zwClS
XNvjxhQSBLgGvk0X7LK4WXv5HFDIvy16CZTp8j7oJy9cCkCYaVxkRPZE8UbEHepMKbZhrOVcBgMt
53C8aLdYsR+SfktWzri1rgnuT8U63/2hiSPZ82LBQC6SndyoRO1Hls/WPOpRTWbEPv8UPpQzD0/+
sFyc0ohfqT6gbBsRXh+o4PeG0aEFzqM1xU31Dr1zCceuvCVchADztLnYuJ+VqkLDT0+JjGyXlFck
eF+q3SjgYXK5wkbnflYCaRnbv9CWQmCRogG073OAYoooL+A9+GWUvomf7UZ+e6YhXaZ/YJ5SQPUF
pDT1R/OIg7irx7K8+zaunVmywoB7EXqDqaBRLTPnOrZN69EIaUuNDQLkopikpaPEevo0KujdyRXb
yFJZCBzJZqSUuMuCHNpi2pJr7Vg3US2qlczoZxY4n+nV+7l2XLKQy5tFlK+YAumCGHB7GIoK5U39
Q9J6gXVRep0qgBysf7psz7yeloiYesHvZ+sbZPYChGIgHfZ8hgL6Q2EWAsfEzYcdM8u+2Tqnge0m
HgI59opmO6M9c3/rtIXvI5CwK26VBZv2oxAfYnnkkf+MLD8kibyTJrb67SVkHLz3W07fdH46xpuy
U19G0oWlJT9QYULZmbEymnJGlERPTYkc81qluxglkGtuturtjPnGvo5EnPlPD7TiYGHNaujp+wab
zpthPif++HI8AhPOsOO+VIrp+ZJo+OdRPXI3p8d90MilKwc1OuW6Xsg+1a/sB9hi9vdSGtuP4TKm
JTGEmzDs+9twiz0CkRJpt5QKd4IyY/3kkUNeVbmFTkRTRn2ohL8EkNVlIu5fpDVGlC27VRO9kT+n
hZhggwfsgODAoNPT0wgFkL0N0d6cJVXfjbejXG1qjoxIT5TVhT57SL7BRHgaHm1NZ8sEQo5UAo5W
IXw0lv61lnHEk1VQYzGX4MhLHNuki7N0axhkCztgh2ysjnWp9yyIDt4ZWC9ZC0NpVymdfbtomEjD
1CU7f0srwCbgdUrH7NH7qwepVpQ+LyxcD1zCW4/Ax8Pn+eu4pY8ZcPnBPJ2fqD/D8NN47NQ1JQOy
KwTQz9XKygqvnjRBP8Dhf8YiyGJSi4ZrnvcipbxkNW/DOwHydVhruFWA98sXWinAVAevQlQXsmde
pVWxKPrPqk1oDPaiQOvVagXB024DGgDB9ZPeO9lV1CYbw9FQsTS6DnaFm0yvgilznDmUrK94R78n
b6sSBxiGQqThdiUt3fQbMyeyO9HY4DqzNpx3CeYlv1p7Ja+jV8KhSCBgkVHHepM2MWRwce0NDOfj
PjgePVviFhk8m4Cy1t2MhVfz+3A6U/WQbsMqH/EinYJGFozxKUe2yfAfvJoSlImxIhrv9/Zmokl4
IaPDS32tlNOGA9vHbWRajFbHt5VWHf+5iaqGkdNWnd40y48PJiohNEgaaf0j8K6mdKiS/bHz/10R
a5jXO0krzPPMrrWYTJbmM1ZGTcggFelvAeJf8/shm1UwpziS3yAerOvyVu2d4pmFOAVIKs+W8CG9
bVN0rMa/ip+Uq8wGKG7n80jkFhpijRF/13BPW2Zz4OnDiGc5QzxBQSh+n+z/0NZqTG+j4kxr8jmB
duXLLyKb89BXp51CaPgCtPvYTnMWYw6EChRgQQDSxgGPRfvJAX4kiWK7n6MYHsSFFPdst2nbTCY+
bpPefbE5U4tmltG9zgmP55rWHNkdDGYK06oS8MWUxn+LGNyAJAgFehoZr70bs6ASMtSxntIKOJHt
CN+LNExR72g+gF8U4Au8YGAy+O074TNZDjim/ucDy5GqgVaEKYSSij83oT5ZUfSsbqcxPY56GbEL
SEGDfUvUMtBsh57CydY1HqWnedj6PLrlzgyXTDEhzX9ITwpPyCnMLzNjezWv8KKN76/nQJa8XBXE
za3P9bp4x7lntmRRBH1HQ5IWAM/HN4UulcmLAj6oqGh1pARmKKjR7qnkeat/Ran+ezLs/6YZgTE5
UcuRX+R9baJj2W6P55504V2ujzk/99k/FGFR2inqZ7CNt8TD/xwvKJzG1CIHEb8hFMnAeZIagha/
c6WJt1DK4hgnx3H09M8+RgY5pMtpwr1wrLm044KzSkm3wrkdF8PKwAQcmxPFLdOaemTEmVx00KqE
2DMvDLQ8+4vwbMPwUD59hk8QuP5wDlSuBb60NoU6v+s+At7KgRqZEKma9hcyvXHADraffuaXaV+k
Ib9aN8AMtsH32vzeUq60oN1QfT9L3vT1tn9dRYvGrEgBgCrgmf1U4Cy7yS1nBfGPc4GtYwG68S8g
2W5A2Eq9nsypBMlD8fE2qytHhhRvmPHq/br2DAxcB3pS7NoxkFaFpFYtm2+yCit2dpJ0umHvUD70
xwR1LiC/lEGppRHjsBSiLlf+rhGzp6Fdu71o5g1OER1+s0sFsFVZZrR+miEt2+KvsumxSLY1ONDn
ooFJ2uOaA6HNjfOu/XNH3/JP+HDPg3sMhUy+DgH14kYTdxPjfD0xZVvT/nMRi7JHyCT2jLsYIZTT
qxwYXz/zQpc+uEE12m+nwsSTW+hK1eogMPb+z9ilGlIJBtIF1t1a3ObyzSkq4UR3HbZzNEezHPll
ZcknPU4WzgSJG/SjW6JxbTfDG/cboA3VcX22ok+C8xLs+rhmkCwpZaDbXdBSdSl3OHwgCAXKoMOK
aQzjn7PwFxxw+j7bqovzcSP3vLEJHVBr0DPFFI+B6rzpf7Ko101V0g1OWfrneDrRclQBz6+Sr9eg
uK0Hdn/X2X3n6wnECfprYOk4WbkJSQrgI8trKRPwwtC+ecmVx09TPo1yV3rzHXCTPg5paTqHzuAo
z47znj+TR2uZnmnkV70wG4BeLbpmfdy9Zqzzxd+zqor7vqwa1Lke75pR8WPz6AxYMojGOYkE5KTm
pK7SZKpdBsq/SPNs948BMgKX0NWm5WoPjIVQWnp5BgUCj8mWJG96Scu4J/pTZBmkjurotA51BaBE
QwtxwpofObu93TEkGbjG+Op9h8AoUUhRaAvYJ1X+SDklSN+DQW8Yh7SwsFC5BErj6YGyleZcSvV5
1W12KZEHOYqwviK4+SxF6cLzOz9Xy3UgpiuFPt7wHqeL31r8P6j0dsloSB/61jf9qjGttR2V4ifV
7y7F+9JFA2nk6mLKQn8VOVy0xnTwkI0OHJ9OIAtmatEkrxEn3zCn6T41cUFa8QGl/mti8+PsWWLV
SO7Gv0feqIMQB3GMTES/D264uOpdlTMfDuFasrDgafDosQZXuqfRz15VSKB+pkkNtQQVF2/EL5S3
Yj7OChpP2XOaPmnI1Ub91Wqnxm/vCClcLVLbXhk9VaSUdj22Mrp9RyfWGJJ2mIHcHAu03syNAoQV
pwnjpzmo8IPRTP7mYbYMvI4dAD/J6pwpukvOS/Cv47eYGF5H2SmS9HJkMJoXJiy85guk8IyhOLuo
3CUnvM7ARYviVl7MZX0o1rtegxe0WYZrG6dWtbygHqoHzJ/mM0tOqtsVuOx0JjgbeMjALldxGXrL
UWReL9OqM0oqhEzGwuQ+whXrJP4mloImN/aKSI9usbbjpCs56NE645xNiy2ID+sm4I2GKa10kvoW
I8h5QWLiQ0CDjh1zKaQZjVIgKjM/ej7G3O374Z56mU//+8LvKUQ7R3h4oLDewuxEWNEqAfpZuFOl
NILWG5CqZfMeUqXVmhna+KPix2ZvQgw/QMOHKZLZ4O8HOu9j0GqEVXf61QLpvLWYw5AlrCe+Ih02
2kcLJXAYhO09PuE4azQbIeUvW91+o6pbbYM00Ok+9WfKF7d8iEUVvKG3Ky9iT8iGlYFFF1agR9ka
d2I1722ZaB6+HMlwu8XGONXOpgAoDiMvCu2/X8n8HleT7AbkBdEji0qoz0hAUxAy1t4Pncbkb4RN
sT8vjPlBvM8Cxi+zL1cdpcia6wyK7JURMjjwyZLjyktqMEVbJrV5iNiFcB/ME44p3wEZm+CKJFk3
g0vtV4r6F17YyJQkFefl5E1ggzfZPMVoPtiCCFWcWUi2/UAp0raz8llNAVokozWjLZRX2m7ckYuU
hq7FrIjtyP+Zr5qvVYBYTsQeHyjbvKP2FYkexOqON/WootXChDSXGe2hwujXNBS3PhvvTJe/pNHZ
0N2NQOGP4iQOaKSTWXr/kZ41I1EI7ki9kT8484C09VjPjltzlNwm49jS6ESU4WA4/5CR/seeBwdn
SBZwDp5zlMOoulLlsG8vt4cl4GihwwkvRr6jVVlwNphXNto7xX7ZHSA/IUUA9A13ZoN/v6oK7wr4
Pns6SYrQERFcCepVYlexTfIljJwata/Ay6ZW3aTsC+yoZdplK/zPBJzZLEw006Pj2y1KkbxxcHJu
wsCb0v/op+551CjSC5D9eYJA45lYyASlrbQQIU9O0LufeKZy4lYWVg+mP58l6oYnlxN1EIAGkkA8
hf/Jysxk4CYX8jEaNJozACzw1W4u23Dar+QzIf0cCybOvaexwPepN7GdUeYm6EjxIpV0oryK+ogK
SaxrUpFxZGut3JhI1NpHvLj0i1jicvvEcxI/cfHnB1uvNBy3dL1+ZzNt0/ZuKGosNApcAjswpC6+
shziPN3siy92CNm2gLkVY/XZA2CA80IX2nXcH4tjic6rrvrR71Ygs6fUp/YdMVdy2ENfYnVevVVA
USySOJWdLPCLg70GgWRtUAmJ9YhYiHI+VIeIQIphdd6HgOTSUDx0xMx773Gv0/AhN+Mpnt3no9Ky
9VFCJBGFZCHePDviGdMmVork93+GO2s+cuGVftBirPAP41WzM+CP0fqSEtIMKVQWb7FwAU3mrX0Y
IakE4Nt4TMR+WpxSgzSgg0ZDS0RBz56jdC3j3yaN1lhePS8RFczGSM2tzYY5Gd/jYL9OGneaZnWD
YFU+F7yvEtWWmq8XQ1rdXSJ5mIxnsDsmTGuULqMd6JtgYD4cus/1pMTL0B9QmDHyRy3jdvSZRfzx
AL41tvBUnbY3m6taeZ7rLrrsYPsOyXMv2SpBLoxCJi2d58zi8f7OE2glsOuM3sA4J6Kvi5BVDtDi
LzMu70Xcg1tdBeBE9O39SqObmZ7PhFEiFPyimVyjZmSDxuxx6DXR8o2tBGE/EWXwOkoOcRyLsZi7
KCjIDafisThRgKxzHeNwFH4+W6A6JpAdPEKYcnRQv0cnv3gDpvL4iab07L3dtfBF6SUjVAfEyvsa
mjMnywROWfjSN/2xIPbRMXMiSvG+KvI+/BENQHvcW8HUFyigRu9kct+tEk88bnAqUfqoCk0L5f/2
IRqSD2qpwfp/NTtJZyWfiVMVmOJeLAhv3wIE0Hvitb9yPh+Q51stp7BWVCNW0kFVzmJOMgJLyKqH
WHzMujLicCMs1CcVkguocqfC93mYwdHESxghY46HBij1u2BdsO8ZY+faVIEpea+X4glXlV0Qz+BM
RFyy2WKEhCg5ujov9acgHlm7/KeMQwyZAyKYcS+hvxAEzNQuiNgKhvKQw5wbkykAPZSWl2kgs4P2
wekbrYtbh1CHchVBVuZ3NtEWVeqpKU/nuRnZjGpjIzNvofG/viGZKbdXIVfEEitgwyiZTyPDGbBj
zAO2cUZ6PlkrPDNPdQquAwOE1+sej5c6dwTUOxljCoERZKlmjCgrMqfJ+OnuWJfCaJSif+io5HRR
7dlIyX/3fedgp/nsSu17lxG5hL+6udPqBOPYF41H4HOkYp0awrV2axdOU7Yjb/vBgUwol1T3omW3
hB8FunYePJ+l1lNpA+nCN0dH+HZlyNJ3vVpldeJXVON0cB5rx5GBuqYhcfKlJSm/oT4VpF+bbEOv
ODycQ0+wwrnj2h84XAQgiYLcLHeNrG2fU9ceZc1Da/+QBctHEwnnIxOyy8okAbp9OTzr7DqyYOZE
uBkJwAL5SOzZ+aE+Qo0AWnkJyq8F6tAm+WgsmqpFRwI50M/jeZJPoJG6sblFaj+yEebW4mjLUYJ9
/Co8QpAk7UPsTDVHZ80b9CIQWSsksMtTVe2ZgniRkHlkLtOdyTOzTWKNFzEYP1sU8lhByABR3yVp
V6IJ9PnDgHfdYRZuexNmXg5q7gDmXT7MIUbFkIJkH2G6ohZvq8QDjOCuZNfjQLuKlTvF3ndOxb/R
+Kb/POUQIv0GO4a7fvFqOpav46RHg6CYCcvuQmMj9qnieJoy9CAZ0hNXLq7qr1jwPpYvCeSDmrML
q8bJf+mVokPtX0bGKWuCDs+8kv18U4Mn1wwOBIQ+GgWqNBE3cv/9gKRl0TZsl6PlT8Xmx278XmP8
yJiWCfrLfWO3J/Der2QsCRSEDkWZLUWE4h9pBhuMXpz8npmilRv5PYOsHga7CIY/4ANZXDx0FSz+
pQM8cdLaRL/IMCmp5OY9NXF1ln9/5sUD6SSSoL4Vjid0Q+AhcwvliUn1GZBSn0a44CxevKFYlvje
3kMkBraQwQxnzHv/+71p8EisIR/m8IgWlI+jga2mlL/fqeQ29WCohE3Ya7pT0wWVGJVaZdTBES9b
G43bLTv+v8fyXvhNz2G3Q0IioSsmfZCm8482drQQrxffsfFsA8EDPhQTtsGv1s5ayb1rZcowoUIZ
XKninFQ6d8laFYh/pFEigUX5yHV2WZW0vtknLUzo2vw8D6bnk0QA2L1C276BWTDLhmphGOSc+xVl
rTb88lHxn85rlRSVYTRctraDWnJzVRny6nw6LPLyef5tFJoXwHgjgmH5rTVOGyV7XpdWyJJb+vAo
Z0YlzKFBrf+DJCwmx1V4+15nB3xxkmu6FBra4R0KvcDd7xdoBOgtBXgDvQZBgT8aMTeRrSgYEkJz
mbV5/CnXyqGyQEGQgkpcx/oZn6qnXrKvVrvwT3IlC8VwfDDqN1xNryTyJlDBqs5USubAGendNDu/
t33K82ZCW25hikKtok5aRs/VpmSF8O/CWvulRh4Ij9B0/ywb6hs7qi7U2usqCSug1xCaSk5tO1zy
+6eVqJkLKWrsMJxx89Y9i/MK0iMD+rMO3VuL8zIlq5Y7XfEP9FIRa1KQ+2qHjdiM9+GIazkCqB5q
zkLLZW3FzfJNHphad7Aq0irB73Y71X1fMzvZhlajc1VDZbERnEYu+FF2kR+guWvcSJqq1QTNwMr5
iI/ff3sXlMHp1Cyj3eVZvngtUt60tBtdHD3lbVU2QOMgsvcrO1H7Y8ISLZ33mEdIayumc7JK4SlR
Bj4Zw4Yb3jbkO0oD1IbHNtzh5+dJmn2gn0qwn+Zx8rsnshovONA91lOlaKY/3nTklNM/f1rchEnz
gitYl+Hz+la0qHc8mlbPljelKZnsAjzQ26saYFNRsiBjDAlIxqDOyP/b7GiMTLoJFHGFrYS38Tgp
5wE5NOEb3iUsUL9nCHIrY0KVVtU8AS3Oin+pyTpCUFt5u56mnJyvOd5la+C6nDQSD7aJdnGUckx0
iqzclTLfge3TMnIx5oOSoytYwgedZJ5MWQj0OF/QEUYS15ysiByDYRpxE3jIJiSrAA0eZYQs/FKM
vk4x2xkg75K/yDwwBn41vaGSusABgVoZV4b7xNjlYW+c5kuOj6Irp72rO+zX/onhDunJqNP8fjwD
KU16+MWagkL1WZA+esJVXZgzGPpQWru18XEy+E4KPymEQBmBuBy7rIETRfNNJQIwRNFUGp44qski
jlmJrEJ1K0fcHUGvjCulK/x12Ev54sIgL9wn/3A3KSQE5graG+OS9WAObkjh/5DlclKvo47yFznw
ESqCEJoSue/aMTOPH3bXxyiNswXeyz4jBKuf7+/fHuCOrbJdeuz3QgcDsZH4juK/+pnMF6sqZFbn
vRYENzCPlKhmTgt88t9xz1Ec5dUdNDCUO644624fH2QEjY4GHmg25lHlyebGhbQZxAiP4tE/EaT6
fSSbDjdXIIRu/LClaO36OX2TSpYdRyNaw3EyY4eVLvbQ6J6p1i1BlimRg7ntw9vpqfi9NsY7BHlQ
dQiUGkiMeKDNksNmZJN898x2jF8ds8RcIQCEoZGb+2/m4YEbdBdJrPBGwEjsAbTjv05i4QmAXAmC
vgApHmwuLfQjvj3OcF04w1iKkX0hwokale1TdyQTpSvof9MnIVIroNtPHiiyV2xaw2kxzmQEhIa1
lHRK/sEDyOXp5QOuILJs1LH73nYrd3FagMo3p59+69yIGV7aNCUzNasaJcItmAZsJJf14B2KL/eY
d5Lj52wTZJcI9LvNTcLZuBLU0NmRBMO/66ECS7/ST+HkBhs4KZKIkp1Rzzw3JbE582CTCOgsTObf
57MmCBDF0WSD9QcoJnTBzZSheN1dF7QNKeobfXNLA6Sl2bQzeqR77NKMxVjaJoZxCR3duJQUvjTo
wfZ+sVukfZMSCj8W/aknWIXIb9Vvg0TksTJLBqOUOcrb4LKYMBjxGHBrY6kGDbn3D6w2BrKL13QW
cVNVTHRBi6PzEVBuOT0HEzk7OBrDLX7aXUTnoKkiMuQFmd58NTlUe/pBwytFuP16oM3s41r5+MXO
t8Mpfg9CQzhaeC98C8lcFCs6fW2p8vxgOALJZTX7e0IA753LXEf1x66cJKSwzGzq0riRQN7HW7iQ
oOWYfHW5uM4e5x6Uyg3CgQPyuU9Sty0EULG1o5b6nDCJwBnnF0p9ek6DJxjbmUKLsygcPLCGICGo
56o8kLjC0UpdFrJDJ1Pp9Vv9YUD8y9OE0HW9NOyHr6UbBjl5BW1uMiXGd/bmwxOzhAgPl2Qxbmr0
wjrLd/GKPIJ5TaesTj6gIp0SKzv+Xv0Pq4RT0XTHsHL7xw/m44s+RNCk3DRIf+O8YZ4o0a3KQUms
1PAH1dt5melWDxm8Baavm74JUmg1N2H96VcZuu/tprhEIV4pNQtLup0F70NVpjcna0hTXMOcQQ4n
UMwkA79ObKvjIMX18aYqyzdqlpjrrRnOlPc8edLDR+34oLmASdYAFinBGIiFy5wq3iVHJNZpsQZe
+TTl7hKmb6L5j9+9qbcy6Yjn6iglA03nG3JdSw64WaG3HCAfY8VRqY7bwpCOaGz44gLhlTBBu2gE
n8jijY0uXxjYkCCe6SA3Qedrl0xE8gq+1Y7rBFv6SVOdJucXJzN4Qp1qenMFGyow6ywOWjzIWKA1
3d4wQLQSeLGjVcdAXV4YnaURm6cJO1bYsb7iFmROTJoPqZx/Pftj+ubtNIVVomTV/o3fIZ3jY6m0
H4pdz/nx3CHFOBpXb/VV56kQKcJ9uQnNm6VtAOAPXpDHfoldTaIltFWy88H7oRUaRX+Dd4DcBJh+
dlOEuC7ho48bwPI/857Lkw1pffOiYUlZcwDg2Q6LTye8w28q0YWgu9rQAiZ/zjMJwQCmZdhy+baE
xxs/Z++leNVPlkbvMi5XFZpo93ZYEfsft1Ei5x8FEMkqOM17t7M14hQRGQHR/xcAntcKjFHzmGeX
4sOZ1RbejVhRPuvLf0mTbw4xL2m+N3ucBULpS0jfThEkBRcqrRW/W/lbwJoAmFpKQiHmbJ6Ve2P9
eLChF/kG2X/YEhZMaEDmiwkEKSO9AqEHjuRes1kVwyJ8EFLxxoHN1rhgh1Ea55ZfqUxXQ/Bo4C+5
qTKj3T287vHutqMAuaBCyICL01DIqIR6ImNAwI/1DEAjNJWddTDlpqPwh3JVYQyp/mrt+4BHF9JH
x1Ojcy4MGF9piQNkE9B9/KFrPrfPbaQwgs/XLm6cd58Z/ItQSJoslChTImSr55zr4dqx3OOa92H2
+vJdReOTb61Zs4I++AgNJnj6qA+OQ3QvOSHQkw+W+gxBVTbccF2L+bMIK+cm9pnBxlfnixEwbjjK
3cbW3NFhTmyVrlJ3ZyDSotDYx20U0hkaXxRk0GmmhdaUh8k0KuGgA7dr14nd1pysKtLf+/FQjDlh
m9BoSMN2L1GDiRtbSEIF0ck5OgodKzeDVs8TxKG3NKWtQRCMOKtWUV+4r6FMBBcdcDmWmKKI7Xyc
rnwXgTZJeIgiMhZczJWE90isr/4zfe+Y90OpUaN8mpFO+cERdNM7KmnGAvWwrMyj2936lc8L8elM
KmqERTdzvMh5DB79kqSBYRnMxPLKzaWqbWsGXE3PJB3VdrJIiZF/ZCW50XKn98fqC5C6Iy1YgGLH
KFcVGrj7puMjhx87+DfPd0738/+w0Hw2HVE1SBoF8k5IoTFnnBz2mjkxDeDtiI9mN7NJO6doNuVd
SLuhk+344bWD7xB8k0+0TBvicQaDl/AWgv9xsel5KBS0Vevyi65VYadTLbgoUPTQg3Uul4a3WPD9
6+xywxHR6fxKTnI9DHNx9n7cWYijmEHisYzx8qXBiqikY9PN9LJV016iSM2+fm5qbJEFnY1hc6OW
zsH6ECeh2IqsE3AT7Hk2q8k2RF9pa25OE1ZeB8XVp1eo8zSTywUBFpnwedeOcfT8ZiUNzASAcq5l
GDU8IpatRip2pX4IcxjlpFhn8ryVdq9m3PeqdBbyijzLXXszzabFTrfW8rnZZvEJkn0Nq6Fb2a0z
aTrR3i2NC4ND5Pm4h7dFnsFBUqy6iLGrPHuhOyFOmegmgfWPU2GP3Pwgtx4xoFCosywWnlvWfJEA
ggNL49GwhdEc52agi1UPfG7/wAkjkwGdMulwBVbgunmPG/GrU5R7TU7//E6HQX/leDAB8R1UHG5i
jas3Ps0doyTMgZFNxIdvOOe/AAEJIUtB3FOP1u8VkWv6Q05ieYVqJMJbCQr7sifoJ234otzlQilh
0BtiK+ee5Dhn/60FnwaMNLq4nyyBPrYpXprzKFd5S1cEc/juAAPQmCjPsq1Pcx7ctO4VFWiZEA+Q
8z5SMDGDQId0HEZ4D+KYTaCZ8pLlllqMMLT97p5hCtJaJE4vJMwDwoRf8NxKfv3DMc33kKTWcyHx
wteXYDklIRAdKe5U9DjGEqAqBV0oLHtU7p7TrQLkIDGDxaP81gmMxVltnDD6SgAeGNmZATsHhCNL
ic80b6Bngr0mJG9DHhwZIAuXXxQ77EcCXdbIwuuPiVg8fk2MtM+lFgucXQu+Pihz66LASRbABe52
wBYyk0xaTB+Pgd9Vl3vR2YipGYo6i5huoiN8IZS1pEo3HJDi6H5SnWgKZQBhRSpCLYIT7fdI8FWB
VgRtuFhSOvc0ztfkrj7et4r7ml5YImY6rGIV6LrN2rHOGN7YR7v0pi/QBqiSs2hicvwxvC+5yom4
IFTjzHJbVyRwq1rtusF+liLgZdlffPI/l6PcTjVPnyc9PV7X7abkc05s4UNze98wT4BLoGfynW7r
l2AqtmxTPo3HCw4fqT8rq28eOwJ66kknsZVgP+1sQtyRfC4EHzDx+5VJYNejXJ9i7Gs0Kwo1mhk1
2YnA7ZyAisgvhIOxKMmmQFQWPr5zgfJobOr1r226q4zK8AM3mLPNFLTUd6a6cEFjW9KbDTImuRJZ
vE1zgvzjZgyB4ydgoPKBALdgEq3wMwQy+6TxXInjiwsqjggNswW40aVvqUiwo9uOgjPPbrfPGRxH
7/1HA+XSB3MUeFeY9cxIq/rTffL8tXn2oEpqjrW7BXyvejBm1oeysFjBge0I42Xv+KxQr3Gwc4vO
b52ctBqZ3VVcvRthCbPZhL0ppwOv0GYgHShF63xgjGSHxaa+SvXbdD4u+kxSzY0KiL6NiOF/TY1L
idJNAdQ+SfGFLEqO2ZEkLMl4JrzItY+QPZ1SqhkpJhLAzHzgq73Hy/MDl+akp7Hie0cHM32oyy18
K5UuEdczZSBwl9hluqatMhd4X0NjAtd9t7E0IGQOFEmzCDS9izA8hHn62pwhPW7apAlMo14NvMYq
kBWmijBbyX+lgRNTgPodVmrzlc/aNmelv0XXlsZOf3hDLtLm0/NUZYCQX6Eb7ja9uNkdxUQcyAXp
jI+ccrDVLLl9o3p/+P4AI0hqoK2A9s454UNbNpju4izwfvIYV1aEk1AVWGSIqsiR9gyXS5oLOdon
fkGlOoF01czKYUKqC/h7aKgwrQOkJLbcSZ44DLfLOzBTg7hPe3DLzlu9VDOwOILuN0BP0yWGiefD
mUzbLaZ27pE8VGwtQ/oTr3nKTb1SvCAXErJCkBkQh33IP+hoDL8JbfAl2eSKshg+3u1Ws7VmVLT3
sGrD1DDuqLkrhJ0NRhd0t4ne0oBGohC9lGV9Sc+YlxvJsKZRWIlxK4Q01+XmfAzenIHvAjeE6zjq
hFGI4YGBePeG0X4TQMblH8uw6mS5pklAkd5phVm9SYV7IbEioP6oSwCTUhmilQPS8tr3jSvkFldM
AJbJpTDMY9vQg7ROhi+E1k4s/vS9d7xtvRRtKLMPMIGxImYxKzdN8SkDdRtwKBMuliLPslV4YEuV
zNmK9mv1DaCOzEyrMn/MA4nhrsoRVq2r3UEkoIRRAJOsGGncKz8sfbhTKVY+tFIozo2JOSSfI63A
TjnwQiLWOqdE6+MS8FhWxgL8wtZ/XNdk4N74c6gCtlJcOn8E/KIc/8LQaLwoSKdHoEWmtp5wr1TP
Xa2qTM44YnloXQLMvPW8g0sva2zia9MEMZeL5526R964Y25bvEYT6yaM3J+pHOMRknLeTG3cseEP
NwYjuXdFz3GAIBMTcN5ge5xU8IqEmbMQn5EyQM5LA0PHmjpUwRe9dNznwwdimuuooFOadDxlsEJf
+XTwCPfmLlVln4tdNgru8Xn21H/yHUkPSFHy/E3EGVvyrSzGrFAvw26i6SaPGka2Rl6IpatBfnFb
hVLeNTS0pPRDG43DgeAgUUY6ClXv8qHgvhc4xh9xjWS5FxWAsdVt8SrE8wHQ6mE7vnhgizPC6a4X
ZucP2kypZU+Ea8ExcreyeJw0NkjhnNi9TCNQ0OBW/+Dji0bNv3KhYQsMvraulTpS38j64Hufpd26
9oLB513W6Gd9keeQglcczV7QDLd58/E41N95ZWOBufvzTyujQNe2UXE/VHuC8QurhArtJ7xB4MV8
8ywhXK63bHWKDfkc5goLm74KnyfVjZdtcIzYsdUFYKE6APDTRQ35OHYM4/5ikXzQqx8K9ZBBB1OR
QSsbD5O9t2QsbKmxtmwZbS6ovIjv6/EnMToV1viMkYVNeBxskIU4wOR6CARJBR2eOJKsK6c9MYsn
AWdLa6/iPsmyw5+AZHe0/1BYTvqM4wIGyCFN661h54nLcoTjG4Vg4M/Ll7o6ETdFUPAJmf9aYZ6h
Sr0ggjVC3NGl4hdFVv4qRIjbqA9ea2E9UKGvJBhYBkeup31KSScCEzDsEcQ2M6kOusQ+P2dQXa13
Qw4jPuki/Zm+HVkq8NZ/cdsGTv/Jj9jT4O7QL+HNcK+kf8FPSrT4L1nMlWPuMQW+iAwFYEueKAEA
5cPahz0ljT5Afc1iY/PYKuixwz2T0YzXVw/ethWfmbeNGI3rd+NdHjTQuMNPdsXQL8M1ItAuaA8a
EPYeUQEs/er9l6IlybBlxudagXPChN39hTKVeZHGlMaMRyFAVl1VMg0GKyv5ln9YAw1L45UR0CzK
k0ZS4bAD051PZc/nQbefCG4dwvNVNkfRlURUSucZ7rzccQLNAhDRY/Biv7WXXth/kghZkrlll9A5
hPt7XV1mb4R9GGOzmWgwSJmiW4VHXWv2o4uqDCWAN0r4eLHgPBR9w32J/Lq7hiuHVqTTKs8t4r7j
YDgOvnODTZwbhmCTyJ9uAgoIMzvWHielT/w+FPygfu6qD9/6x1EO+79l5Wp40ZCCB1px6LfbIbf2
gJaKmUK0plM1uk8Vcrj/eEO3521pP/ElY/6X4rBoy8EHz0Zw+sDr6lOaXuYRc4FAbSingLokHRQQ
0q/lYWNnh2laAazrNpOZa2sJT9a8bwCpFKDKdDn5VlwN92j5pxSNmmUrYP0CnUSZZOgscveeak0S
bn/5ui6v0tW9tKg5Zd4I/y06a9mxPOVJ1EPRwzPrT5FiTVohzJraxQ4jkzyAWbwdC0C1hqkwnxDo
qHINJOPb1j30uDNYY8jFUDTfB14ieBzASg4PBIrM9gm3J2xyc+5wddyjTxuDEdKycG7ZRnZkf5Eq
zsOoJ0XdWS4p9dMV8Pmsd91Qh3c/O6Ux2dtC7PhgDiKnAqhIJlN6Jey0H/Bf0rhUl+VslZ94EDM5
/SHt6Ae4zC/E9SJLgg5hHkwfFKTUDTaCi3l0BA2fCfhxG29kHf+PxiUoeoDx563PES7y9oerHemV
znI0veFfxVs26AhCqBmN/TY784Z0bdxZvV+nOwYTPWMhNMKmg/yCIKwYYvi37O4+zUDzUvgHdpwE
mVue0sgxjppK8D/CPpBdDUS5qJzHRHnJkVhn1KkErgjLPoIxC6xJzYfTYaB6AnkwEHvyuCM2X1i1
kWd9X7aevtfK1moo2xItFELaoBguV+IqPM9mLyElrC4wXeIo1/gybPPWGF0ZtXScN3fTo0SIvZw2
f9Hie9KNhOLnFYNqq2Zdb/n5qd2ocnXpZOLwDh8CkJcf2t1OLcpwlsjPL8zJjQOdTD5tPWnSwRuh
Udq7za7X1k7qWnnbIvxGkjPuUm5J3rKH6bMDW9wdK7jmmg3cQq9efPNjPS8XQOM24VEs3XhyYH4J
TwHuZrtFLpT7SfRu11UtUbbugTbQKVY6sJny200RhqDDBQNtvUl0nfHvqcyTQ+p6LnyY6rKU/5iM
Qe0i8LPkGw9sMz7yNuMkBrYpHMA6wM5mMVW1G03xRF3j5VUum+cw3sNIN1PjdVwzL96emfRVFaiB
ulriQnEAYXYct4VSwXQjHYc7CS4Ya3vrRnKmAGA9NNU68LYm2RRSC7MnEWpVPolR0XmMFaQQlnu1
RTUCHJU2Ob2MnJclwiJnfDnrmk2DTqQ7jHLnOsq1FkAeF/4AtK2gD42EBY9pysXd6Unta4SJn2XW
INZ6KKjLilEZdwu5zgSU/SjYltU7gHO6hijkkN/Vi90FsfYVeDhH6ZFRosKL5CnaeTVOQmAwG0GY
ft0sX7fs9c4ClzzbQ9fXydeq7dfuz8ICoywnrSk0HuNCM+ukusW+u3MfVkjUz5OCjEzsbDoke73J
aT9VxICTfE/gnLFTbDvFMYq84RFnZ5bZuVOICp20xsZebJOMM8viQ+OrRitRxLissesMYqQYbi9f
H3FSKMMbiNcchhzMsEqen13rVsG1Jn0t3OEr3uZWJbHiV19/lcwQeBuCZ/UL+yW1SNCiAIuxJ3n8
rUMo0P6BJ6K/xP72Hmu1ol8KykQQeLPFcR5PV0o6BESwOE+SBszdtBz6FTrDfNrnV48tKYlfG1xv
1dRIKrzTr2i4x5UG5rCiwqCAU7CKFtulegrH5AAsiZXtKBz+7R5NX7b/K9DVGwnH7MSpYmLpSj3K
eMwcXT7qfYOEdC2c5cf3+vbCSDASKuzi0p/kSucH1Gm6i0ge/BIlEM6X90ViqO+9jat3mDNPLk02
W2uF1X4RLclqNJYk3AHn1rOcScZl2LxfdNH43Y3LrZvjyGUBoY52LfPK5+5UYEvKma9FZvICwJ30
GhDsXrUOy4eTsjtoV7A9ppcJ81qDj+wmoMvSau8W2t4iwIPc2bINRiRmIz8gveZCgsErI7m1wdw4
PcK2NLT9zOwSawVQJpu4fchEtFsxd6j9O6YxfIQyZPLuuyv+BLYstTGwHmXDMAdzfzFzbrqzCjDq
SpN1fmmpEANC1h920QqPGguA2RR+k1zRhiu43XlO8tG5XvmAIxjXbg28SQuauetKJei8e1TAUfLG
lQemDKlvGjXbFRErHLrBuXsQvsMKEsb+VhKIb6acmDuZ/mP2IRMHvIKOlVP9wUS/I/wHVonwy15p
pboO2wpDC8fYYv+oJ+E7dN7K6PUWGzEW+h3S4pj+JWT5V9ln5wF6vAcso7ttLxQixNLPOBftjuUd
8hZw51EioFbj3z3VrQBw+jT4Lyb9hFoneT6yDwPpGk5zw32IvNtNMzrgWQrT4zSL1E5ILkNdNIhx
qqpKnsHVWRn0gNiRkrqp9dnEpwU1DzM2BX7lEv3oar+QVq12xqLn2R6LKTztLPVy4PTGYjtWFKyY
agJat4XyAtwp0xGnhSk6riAt9hgEpP1uMOchhE6vTEb3gPcUEXfOWCDGaIn6LbPvuVF0x8P/HjlP
bqRXKTUf1/uVXWtyuocWTwG7KHj+OzHII35rKrJJ7VlXimogpsykWr3JsmMqj8KZw+m2YhoVfUBW
zXPIVgGqNba9MZgsv+Ug82SU7KUhNmJ/1iwbvIFvL6hHVn+uYowTeyHd5cIaEGNGNFzBZdDMPhmG
bn5cbmmBEeLmj5ahRjmt3QbxYg6mICSnOLckM1jwF5oBrwXccCkAYtKl3JoV9/nzrIaac2gkF4WQ
07h9/UwQtRYz1/1LAsoRTsdrLA/HmCBisUrsDA9/cvYwgYl71HHGno34YvRRsJKQgwYh9xok9601
DTghViyU6pN48m0Z1ZEK7KzzABTzWwF8s2QMwG/NCVohpkQOUtZtkZi6EuS/MYRPF1glPNXs3Hg8
PxqcyCLoZa8ef60gIbyLW7V97jFVrj7KDyZ+o1mBVLtlWHdWQad/F1R+6kBgysBWDxnPShKN0bnu
IZhkoh1vtg4hx9/Gw2bt/1bmBLpmc39UT4UhC6ztEgo0ETaCEO7rV1++UrIMZnEZZ0fYKnPL9EU3
Pw50PtO7rLs5Eqj7vAnT5VcU+K3v7ImmMrAnr3Fmu8tFD/ZreOK678b35TizmovZR5PuuWIbXvK3
iuAnUSKj1uTVke+UgJZplE8ZdIOPJMLnVb5iXo7BV0QtPopGxv+exXzDmcuniKX/3CuHWaV4/wXG
BP5CIu1NHG0MNUSp7QnAI1TYW8DgWvvWniMl2NmgmZ4tCBJLMJOiBbGigVaBtEx8ZQtcMjUcTugQ
8mDyXdgrUcJaDDSZ5ebiOWprZd3xACsyXq/DqGWqUB0msm2zMAYivD08WU2gtYtzyQpYiSW6csFe
DMmti5a2PRJLcqX2gog7NWnMuo8kxsdaKaxUweuQZtPOOqbUQy/OM8H9iVGRPXhYd1yXFvhEIztA
GFPmMXRDzmpnyd1PAdNw5X6OqFxqWiJn5WKkpWhvnRIJoCzljDheNmU92g5jBHHhZTXM0d0ZPEOd
mrC78JFdeGkciipP8LPxAKuSlgayrzvLUppZUPkBn5V/DyY7n5HT3PqUnuT+wzQrsgbL+egIiC+H
egPhqHN6MOSU9bTMhYf+5PuFEgKu245UY3axD0dLr649kzsL2Uw/J6ExAw6S/7yJASEdd90jiQ5o
eq5oiOBvkJMDfaaNR7rHAUEMTdhFnZiYDMR/TkN1yhRVwmjRQt+8GvsDFr9LF4uKUH0+6tPn3Fkm
qF9qxChtxuAoAaMc9KqQAg461VUKvKLMWG0QsPxbPA45/4fvBpOwOdJh5FdbIbK3Z92HMDLgZN08
01ooWQCgWDEidaTYlYkKGBMLaZy/KMHIar7LGFfiSyIeGjkvcfnLYoiomT3kyxpiKQHPJTfU5+k9
D4k9kwfQ1ncxxJg4V5rL8BN55wjH8feCR28rGOfw3BMWOHWCLUxZSIEdcZR+CdainxBzwPijsyDL
eQF0xh6/E98gATEEBu9HDzX+aA2bUrF+ChjHVOqIg6rO1Uc/PYVDQOrUG5sLddRR5Z8fkyweEf3h
2Yyrl68149Wg4j2ZU0KPQIPyWH5E2VzEpCBUTRsnFM3SfaveweUte0E4uF4c78S02XiMcJ18DAKW
sbl0WAxohT6aROuoaCFVPe/URrC5E6PktNiTwlfuJa22qYYNYaKUeHc0ZDzyX1Z+PUOV7IyWygYZ
OCLWT27Gov9+c67jkRJjQ6aM8lqxNT1sU8FX2lmVhnMPhnEbmQH33MkfuSFJeZYqF7Lj2VpamieR
rBlHfGtj+5S30wt1NFae2CWZqeeLKlNXytUrYUujC4XW4lZU56UD4PRlAosntO1j4qHSSBppqqDF
sEvDkgmat7QKk2CgtsxLBdsoGocD9Ew3GQbvi293TNzYIIxDQWXmCL4D9T794o68zp/QWUEj1YI+
IUiKU4R6wOzBe8LGVCdX4/ulnpkaBG4t/gDiC1Rc1eoEE9Aj5/Ab3WYm48OFIKId2k7ew5f3ymyh
4fg3GhCvt3Pgx6KsDYLsG2tPFHchTMizhlWZ4eVUSKWxxEmOnPUrtCJKcFbfvPFE6/jBkDbdaV++
yaZ3pIVtsyeyz0de1WnAf1UvgtYsVU3kNhjolBkEFjxvWUbhi4Yf9NGqFSgRX42/ToDS8AAQBPne
ROsEcDEqHfx+9/Cxb3FNZ0r9ozQ/zwdiGWfsjnBgmtm6C9sTVm5aqculVz8cv+Zsy1+yYXU362rm
OChH6TsOfbpXfXUvPCQIqhwDWMDVslHvBi8+PBVNIpGk8O/NlhMR/AD9pOkSBBuEXxp1Sj7bdLu4
MtgoUtlZuntRgJT6XWyuSLGSpgyULaydrA2pZPHMmOyWKPFCeEv7AvryM2nqo/VsNYWPPHfHh3hJ
4W1bfWLfyZgPlDFfMk0o6bNXdoSA2NTKYetFtXKNAP2ygGJf+LjcMjYBDcwA8K+lerB8bm4H6B5Q
XYbgnE7HcryeueS0RmIV0x2ZPYphqU3FgI+zxaDACW4FRMCTCJLVDn80rdDdjXllMiYsTGKf1N6v
OE91fS4vpJt13DU46MIgg0ep6yXndp90CrtrXyz9L/CL87+uK4nno4prjMemjDnE+E03Gnf+Tc3q
/nggku47DQGpfvYY2jP3cv+GD/qacorqRbhnZ+oM7oHEEFTy01tqLQdGzgyHPW1/OoZIs5TQz0Kt
uF8dcSf21zIxZRYPt94bmM4FKjfOlKOnr5gLzsHONA3i0uAG5TR1sTlHOWmnlX8rUSXwVswKu3/U
kz77q349grTat+vIrFvN7mLrVIzqBLO+Ri/4EY63wgKWzCHNVMcFXv46YEK1mczzPngXf373Evh1
bwIBY+u6mCCr+rnTi9IKuI6oaaaM2j5IwHRYCH2estfF2JYOKCtZgDa0cv31J/pb/2ukSzvOiuq9
JVhgDtkDR1M3emVCYRgyiva/EUDfN/l6NMT25GP1dQwbz5YMDN83CzjTHI0S2EE6/RayJt6Ko9M5
Xa3ZuD82bMGBZxSgTqsakX62IsA6q035O/aKTu+6ZtaRJEt9ZUEZP3IaWuNWNCgkPyr6VhrA7bRJ
i6Lh7cR149qobe7zEofbwZl8G0ASvHe0ZaeIHxw9gHEo1QE3eQPPY8SVsj80U8jkc9jCS5hUeGnX
FhtPsR2t25XRQcYQj2UnVA36cBfcNIzn43VZBsffhMBYtyquhBp8P1GUz8whEjxKLKerpkGVEu/R
1y9vqwYmGBQh9nbguzCyFQW/8l6P6k2lkQxcoIhCtQWRZ4d2aN1JVMYUxihz+EhfNbz/7zgMwPvj
uDQajJE9icga6owhl8IgPjkMZeYi0G2ALZ7PEPE8M8EY05LixmAfGp9NqknBNUSXW5ntkeseFAdG
OHSoj8rACBEYhpzjoTcc+9wqijK0oBX8LqogYsFR6ZKLc3kCQpNgIFk2KeE7dKmgMCgGjbedm82x
rBE+dntK43AwMZmP3H+gkDW/XXh0u/TTzB5tEVhokfdJnybtXhJjRQs7xATIn8tP/puNFltS4/f7
y2gCL2YFuBL/BU25HY6GKjzkFLJheW8picoV0JxnjZ84QF6ZxCoPBR1yQG/XTWptdYs/XeXo3CkU
ireBcPd8SupjO53YCE0/0WnAkU5mwK1VDbmGcrG3uu3Z2DaThEX6ZgJLLEBMZxka2nN6XHm4VF90
s33DxPGCAeHcT/xuFLzCfcKuWUK3S48Pa25tX85ga3PCsUdN1VjsWxFH1HRdf+taZDEFBtm4X4fj
mSotqTuoiGtbOjih9ex59P8AFX5jVllQxC4MOWqE6EekpVqAjwFp9akz85cSe/dqn+ctHuOy96gc
huA/xDuaqbrNOsOJ6plte4tyVh8R7fLRuuoUqSp5FjjHg/DKNXEAnYvw1s4mr/KnvI08i/MOiAfI
KYDMJZ+kigqFLr+Axh3DRSjyVRhzyazOnheaBDbG2vD0k8wzbel8P1ifTeMb2cbAGEJHLAJkqSP5
e2a9KvAVfiMbmHVKanEioonWZWnHevoNMSHdQxMyAtggKg3CqxCwEIB5crHKmcQno/kLeOclD6vX
5QLQk2uxTuTOpOfHUv1oNUHy7lxFRVj9MkmWG7wKrrsxfx/hkPDcfQs26QcSKihaocobGew3aChs
1kRsoA3tXokzmhYPW/mm4w6sb8ug35OzK824FNVUYW/c0z+LhXuivs7PcWWOXOjVCri27V/A0VF1
ZXTB+BNttSQoaxAwJtdNSSNnpPuE8qjPFz7n/8qsoThrDVtk5bIIFEtXABSkOdnOuE43oVfhbpGS
md6GoHMiqI5CYv+TLVMRoM2i9V4s4Rm9hxTRT2+BGGpJzT+dzygrpJA4LgzKepYEAnbPYCvxLFin
sDq+XJJ22SwL7y/pL8nCBuVrKWzeqM3rohaGUdUeZKGY61e9p9sYMHnfjhHt/9o0hFYqFhFVXZXw
te9vDvaMQCBFF6V0cN1Q3XFvMEKb07f/4uQ+j8PChcxXOIHMtXs42rcW0aFBHw0owDdHLMWcVn58
tSPr/RfCplCJN04wCCuXrCSxLhS0iVrtWTA3e9upnMKUrqIrKePw+wZo39eK0VYldt3/UYXpG58Z
8kVuKgxXc0++HIcdeCYyH7Ve10HFGXxl/C6+qVbdv94rm6xUzZV3micjDP53jQJXd2qvNYWH39PQ
Ifj2B1ytlGVE8UaSk5EOF0ufLuT2v+xfWH1WFcAQ372z3ScqJolxIpRIF6aJX4ojCFoLRbJojkAT
RLyDBCLnwoZEmXfLjQ53VST32O9vvwCVNytScWfxbtk5ufqh9YD8CPm4s35B5e5pF2n7p8mmoLvi
Z0pMQy+N7j2r+eE2dKQKzCyX6Aa9MOfV7++jXhat8jKXiTY1u7kxoyxq/LIMR0c3MlW8Bk6CCt0W
lMnVnJ9ZWAHqVk6PMmBb+U8Xg6RT12SNFQTla6s38V93/wIPblxQZh5uKt0puNSrS83T1cRdj38r
v89MuTLOCPqjWL0fu7vKPdIcuVi32YXvoS7u0mEYPp9bhFyKG4iDXTWyeJVHReT8SP1u5CjS4yFM
u48L4hrPGiOMh5YYuunetGlnzub1CfBPR4Hr7SdkhQKkym4tKjmunCGWRpT/SBBNcuwiH+N2SrL7
JtW/j2VwFcsCthgd8HQhtWZLxpLAZ5qDetiEYUWWL6+BqoGo1i8AZWe7m81Ldo+BuVK9IwG/aTTR
Ym7f0IezaZb8Chs9OkJESbM5QRtQk5+kxmuH26DtjaEH8pTTdnUTPDJcxiK32zpiYOiSJsn3uWYF
7plrOQt/yAvRRJbtPu0MMDqiUymGVw2bVHN8NM2VJ58uMfSO5g==
`protect end_protected
