`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DzhYMRp1NqtOyVtIw3kXGYP9uqAESY8bA+OANz4RLsx2Xg/WPZbI7i/HHP4wh2vTbzVCdPuwP72w
t6bWCg1AHw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A4kKK+cmn9Op/7DJQ5eJP0xjhTaqTw0c7l+VooxIBmTQHbezHQsh33vvPcHH8CDja1I2+lKrOst2
0tFXbGTJOcQixqpG72bT1KHcpvGrGyUiDShkkpqm/hPk7W1HtHi2wua7nnHJPbtOpjy3ENFIrcJg
BK+AzrGl8PriZqlvVNg=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mGlTtp4EdlCAIaE9lGjzEjtQBOuQaug6AmtpD/mclDWgEra/jzWgu+e1KMcFuqWf2KpKraIMeiQx
KnNil2NGF9YOYVgkkX492ZTmSxK1QLO9p32dmdkfnGmZ0m2EkZED2YD1CxCeulJx/eQqXUs8i05V
/kf3+fecC1rxDzhkGDQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y2GAEn1epY6qhtj4xKTWZc+3CgGhWbqa44iYBbhYi0GK+6lBmQzSBzyk4k8y8gabTj+fTHjGDml7
Yjb7DjoK0BVA3Grm48p4i6z7jZOF/zllwZYDdQp1D8N84V/hmeHsD82jQ4BzvZyldDOoRJu2aPH6
69xtISwD9YYgkR/Epi99cDXY1hofXoW3I+I51rO4pPWHcu8eo3iI1EtZOmGDE/bO+GUUDc8WA4Z/
Gsz3ae5xEeQFFk3rU7fkRKvgiCwFbCX9BlvNulRnSW0UmqqD1XpWjX2fdUkfbVjKZbtUi3Cmm1HZ
vMa71MUrfeM+hwgHjM3+PG33RJJWLeCq2MWlmg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DvX7eyURz75elY+t3pktyJgsE/M5W2ZfMp/EOoCASciQ/kaPgU7xInJfg+WcGBBbu0k3LTkKA4aA
XW7FTeXNMBRppOiQMUFmoVLTGrHewjrX0e+WFtXdj/Llh/qXcrW+7MlmGu79oGL/Vu/LOz4rJOez
veO8zuv3g/boLnUDn1KTRmamqKIIHjmYxKY1qUI5r0J/ke2+rnKYReibk8DM5lrJypTPFICjbzcC
c/01Oxz65dicTiB/yrLzSddtjJLILFqh+k6XemD0pbY7c0tA0rhLnR5F6gn+iaK0SKeCawlqcPbN
s+gNs76TgGR9puGLJKUjnu20DhxFSiUpNSUgLA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T46MqxRu+HMzZTF0BgfAkwuUC8ZkbSy7auCUVzMxZ6DddzZ6FL0VfteNDuGoZkYvD0Ng93xbYEyd
EqHRcXMdtmlPmhgHYcuTU2WJknUa4FuDV+8FIKQiEuEhvxqYlxUPxcDPnwPpHL+eJlHLpUisyqBn
sZpJOLI9ZgavLWw4LvkV9UGR51BLJK31jsHwUBYKhPS6vfDr3wdyfYYjXbr+HlHgRVxkJMEqrWyN
AmxJxasSVPs+y393pesHnrFoG0uu33W97QEsjsoKgo9TvjJuDJXdEqAUG6mhCh3uYUh6a5i+R1Xk
g0oBOrdNmLCETunoopZbcAB9DX3pgq7Kym9qRQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
HmxeoQzMMFFEbGyeZmDz6KPu6pxGlct7O56fCbjPEJ6jsjxvryYF9b/XLKy00fbJMBknP2/7XVFa
Z2kAdgqZZz8ZJQ9u2ildkTwwF/YEvnswUCMtk6fSlHpLvG6lOsLh1Qo2r66W6iWKYzECyvJGmgxW
m2KrKGfp1WGyKmBsE7+NNfH+NlQFmKzbaee6S9px43Wfm9HsNRrTtOTSbfjXOpjOvutWE1d6VKqh
siVYje8y+6Q8ZlnGcZLBEJZpLwQTC6wAvCsOpxdWXqFnRZbq+e17wCJGq8rbTZ82+MDAxfz8hSy2
CN0+CIeOB05zZDGQPhfteIQ2oNJE3c6U9mSAdj5nra0r/M2wlAt/QqISdZuDnRybvO+2QnclJ/SX
xrYKvm2I99hLaZfYciLBAboIFAFuLtq+4lyeZNFyZXMS7NTlhG9SOoITu8462JEDmp8F7Rr6cBqY
z6cATeyLO7GGVhhYNIuH0SfOWc5yk+tcZ6/g9eLJjmo7HtbNkvV9gYA6vgDh3KK2Ogndisi+1pqX
zkQ/vyrHnYwnqwqltg0iLsTXx6flHkyzccAy4mzFK3qE95nCYioSTEwmCszRQGYVqUfPNag2PvSl
njNqLTIlWvRyKkfDR85OtuAobTn+xHq9Tt0Z2S+ONLv6GniGxXRHnqNYs4oWCBM59WpaHf4D19ZW
pFQys+tZLFg3mBBiRZNdD8sVbYIT06Mbc5V12wbLXFsFqnPBgAZksCC68W93PavXbPo5Jy4mB5yS
NfILZpefoOWDvaWVroEzMfJxeD6Cx/CDkAIgJQIKXsBv5TkkFmY1mpA9DqPaJB9y3BbVENZz0iMH
CK4OdgSgku9qFza4XVujScdByYDWG7b+UHA+U9Gy6YPxlyk9a1KN5UAt+8dC629mKNxUdvZq7fjr
wxc1hbu/cQOqIPfkxJqU/GE4Y03FJcmXcPso/TZLEaukuTqgw8BkFcSpCB7prxeWX6Ptsi7KHH9w
q24w0lEHNdD94GK3jc/BrD6e3gAIPZ04htqhg74kdSMEe+/veLIO25+uJC9Kd0kdWscvFc14bVDA
PEcny6w0DYC06fSCxpz4NWAsBeha9y92SdR8OPkVeldPZFrqJ6FI6j5lO5iy+afN2tegCCxg4hzr
mErSRxrleoClCLE0uQ12VKv7cxPHwCT30gjyinlvIkMaAM0qg4zwmTTw/7oAkT4L9qJR9AhFVMwM
UR7aTVfCoi5p4OynAsykR5STVbrYkaImnnIGPbNt/J6BhwUe7cd/ieIA4o7Ovvs3la5jV2VGn+uE
fTzzPovPIUN7tpWqz7mWuseFKTgZiNTCriz9YNZArouUv7UKx1nvxNrZyJtX+WaM2wojmk3W5rdA
hSovN8vtXYXvLH5maXbk9fdF5u6nzj4fl9cABW4CaD8Ird+fP5/oP8c3oFFkJrLk2+gUt7Rpo5Qw
B4aZGk4xeF3dDdhzDAVotkAQy/0TINz0rMScN09ItAN03qbRgy5jBDzlttGa0IvZFxMjOSvYWMMD
01tStBLBp5IqVv3rqiiQ+EGKQxRuUZ6sF/eqoBw+OPf4aonF3a7nqwmV1vtQwkqzYPIT8gjySLGD
g/U9cFs22xbI9yfE2idm5bAwodHv24WvcP99ImccIgrtYe1iobQVWLgxRBnVPTOJugpNVGgCuACn
0YsC6mCkowt5IdENrGduUpylxuQtXzWnb2+7fTnXM3jqxXsY7dGWK4qJiu/TbrnFmLiRCFRLOIXr
UCJYdq8DsUrBJoJ68XhaabKZHey6lE1fJjYsMQXOWg34E36m/4VV9+t6wnUOOGqh3GjRQdrxm6+f
tDbNgo8IyWJQ89TCZTJ8xn5GqCfDyi7RwsWuV3GyLyghaHK4qNCgZHj1dMYdTJ7XxRzki6McX5eD
ZjxgHg6ezHX+6Zj1ZJEM6n7dldjNUlViIbK/Nnusb7n8bvgh9/CUWgsYVEic/V1cxPOC5jr2lPLO
7IeazNPqA4/zRDT2Ti2pMRvpZSe9ybIGgzgtu5X8MBFntPaXieL6H8LA45bIAp658QpL7rTlosqj
jtQj+Vyz3hHo4TU0wNhF8RHXG+UVVPJ4gUZTPMWadFSCL1tCupRox/InS6lFVywhtaRaigOqvR3v
Q98+8eoe8hmVgbs2ieI07yCkIiRLK44USqx2XX3a5cxdtmoxoh9jt0ey4Ekg+KAXsnPkDE1SXXCP
ddtBPtoAObHBiiIonqk9o+Sw/DCahpXwCEj1kJI3YAjKTcLBJfDrw7bfiBYKn31fkYVO5uXaEgbD
JMtnYRiaOr/Vt0uoxpJs9GVDrE2i+6+pNo2cjKMH99WVKHzozzhVqGUIJnFEeRCrtZB1BD+yMqZ4
df+sU+Bp8Xg6xhNPA4wQ0rJFK0ivpO6bdufg3bxf0aJQPHJJFyw8U2Re7Y1QczRZxy43GwRiZ04Q
fJ3U9NH2dV5iSqXwBAptpLlPahjwzirvIXV83aGS3UdjRvibEuxNkyDQqFeXQFwLPCzXC6HgBKRK
dMi00iYLsFlFezmZSzvOTXXaeE9ubgVM/m6XVieW4FPufnb4Gk+wAqku3VONy/ww8wULreyZhLA3
31hmCg26tGjOvnTVzzQ5r0dKTBJat3z28uObTMyCUHaQW8xB5LHeBaGFHbMm4b6+ZWFrrHSsIxeg
hZO5YnUcwSRqNIemJjyoY9U1bFyAtY4KOX5kH8eBTw5Kc5H6igHMaeO2b1xXiKFr8TcOWzDnrB8B
SCuBI2VQchPqje3Dt0c+C9vltAM9dap1w7Kr2oeXc8La7WxaNxvp/l/i4CuEBINiKiiNjUSqVGJS
SgmdHA+H9N4u96D46e2JH4NycCKkGv4EX7NBF1A/+xVtmJsSLmXo3YWCYl0G4mwJ+6W+3EByavHM
6tWGpudCwgO5xXXGbm124eSbJaJshek0mT0UbG4ZyTqRrx2DbtRguCY543zwU6DEWkfcxfilNKkk
eWCVDPdD/C5dcuPi4kJtWigReig5q/Ly37d4arF9Nt16HxPbbqCTTTKhydSm8nd4IG4XmdqNavj1
kSvVf+qNJj6yROiJyyUdsVm00MdCg6ZpyqX/oXHMP+7JyJxkbQN2RdI/NJr6jqD5xAxhrDz+W1qw
0TcmIgJs5xspubXND8pNlKRBvWqBVUt90LjdqLxBGMj7q+XjLCTdGr4+yOw88ZtW5Yw5Zv1dzYAX
m339rmddbCFsodXCYpe6b/EzPQKXnod0aAX5xdJhvWT2IBbJBX1NjtByE19N8F+9fDF0h4rGhVpl
3fBak97JiexBo0vTnW3e74YmiFKoMdt8ZRCtoc2rm87b59OdkP7XOCTT4MQaCyYUq2pCG5RHrXP9
1LYhuZfYQ/YYuMWHA5UOKBjrtPkki+x7HS0h4yUDMizj2IR6OHMpYU5S/PCF+529QWXEroObDvjW
qtpDvIv9Q8cmLby2G6ptKPH/WQrEEkAxPCqOKGZGJGVfK+m2Yc5/lhuVcXCc0K4MID/QUagfHKpn
X2FNuKNxmgXM7Qj47SLR0jhvouRHarBnuCxbgYG3Zo+XjBn6dd8WiAFzQgYwviDnc65GSTrdPN9G
b9U++rF74eKtmd1AnqSW2IZ4j+MbhAc2GFWCRd8ksKEskWvsEjYzG7wYsr48A1qgk022lUWyvBlk
UdVrzFIRphUfcpsYtk5fKaW5B7glXU0Q6WiCIpDARULzMyzm1myLUBPPe1dKjPipzvpPe7hkD/M8
qtXZ4+O94J0zcB5IWZnrCs1EPanT7cYUF/ij/FFDDc1SRF8H0RwBgE5kFoMdUT3NPl/BBWM5GpUw
5K234OYtkCZ8y6ShKTLADUSDAKD5541M6UBnoGN6io/hs9pJ6m8o/tjPzltHNt8lFetX+GWe96rD
fP0mwwK8RfGZc4LRGbI3TlFpjx1NTRjLG93pcDUowh/TBYtV6UlLS53OLlQH3bpV4zcen8nk+VWZ
OTRXDKmv0KfsnJ52LAR2K7Gtb0yR4mojIKDigxDSuNHuztwQeb8XVIkP/6n1Pt09HNn5yFkr8WL8
4L6CFe1TzfKfejCHzlTQdMlgCGrhVRqbapfT5/OBdm/ve5Bu1KQl76ONV8twNnUe9VR+uX8UqVg6
o+OKeIML0VYmMZ7dPcK5EB8CXvd7dyGcCV2rGeBF+oQeUyOM49aVQifw5PAFKIGgNU93gz5ILCqn
jf63T11NNr3jFWT5/GAQ40qsFWBp1VzeFPHcCjb71D1YjPVoEP104ouH0MGfPOpB1MHV5xHapUGS
/HpJ/L003Ymr0Bj0DGESCOSpoAlsZE6RpGa4OtQInaSLrROFd6JQMRSwIZGKYP3WJn2kXxJnrbKW
gQQUsPa7tGVOjz3IptRFPumKdBtsgiJDdC/17oVMJgAsGlEaO+ha4fHKyxrdhyIjWdCHENl+mxLg
4PCYoI1GUyit7a/9/hvLhZQZq4chfCjE1tT/DhExmvOw6zqMHokEA8iKb1hMA8i4vGuXi00avBKu
TMHjKStRQx+8hlA6e8MDH1LjCKUyjQFdbQExHu8DmQKH3G3Op73npYU7bUMIekpK/vO72zHZK6EO
2rapXm8E8Fr6IVHA+CdPckyNl1YH5YZ+V0+sbaJMrdp0Pj5+pBQ8S5I+A6V7NSXESY7+9vkkyurZ
7jLf7ATGpze1faAk0x3QKel4J/GmMmWEbGAt8YFOQ+QfUH2/Vx5lTOZS8ePGVll8HCsLfpJnNdP6
npTlGKaoBjz34YKuXqY0zxx85Cnvdyc/rGKmdRoy2xxPe8YrCAIP0pj64HD9SR2nZaOP+ZLSFsl9
9Yt8ko/CZ44aeED17ikplH2jlFdtVaTB8VdM1SAL2ZGGfxA5v3mEJpoHJn3lWiUE1VotnYt4FZ2l
53cDY1bstBIwBQ6wn7+ICWQfrcZ41JUooKayqYUehNT+8n7qDe6EYfrJf0lfYKi+/tG1pHUzm854
6/k89rqKMluCFKN3lau2cwuErSozKErd5OWa/bjATtenI4EIHf6VeLdxCX/ZTVeHWA63UOVUpzJC
27zXDgB9cWSIzGgpu8612brVWuy0dHmnJkW/uiZUCPFrxS42vZEZVKL9wTtZjgNTjl2NA+sYovKU
sv30KEkeBoex/dNJP3wxRLyKyG5v3mjMZhqIvwQ6KivSm1pRBxkqATOb+ajjgMu5zX+Cduna0Jy4
TNr+zFd1WWGYISq8xKP852UDARAooGDl9opNOsTUhiQvsWmoZeyREA8l8kcvLX9h5fsOmCsnyC7C
2cIdNVUe61yxguKmT0Yw7g8t54FHrgGpxt2IBvh4KnKCUoHDymkL/CCjY5a+T6xKCpatCdnnuZCY
uILUXVIsM51b/mG23MvDyjWac7c5cbGLStbli8xij93N86XFyQW1Z2dEblMWBO8CbhSdQcrRxDLH
WCy86UzcIxLUKNztwdLwru7KY0kJ/flEKlfIxE8dAVTG+xISnIp3+Wr6Iqsw+/Sq3g4Dnltv/iwi
R0ZBHtFfOE1mNQe003SHoRyOeIB4ODUc3S6oMb/JiNQetmm8Vz4VPhvGcFwhWeV/2JGhQt6oU8UC
qcPQx8GAMw+QQlCAM1OBQKyqApVUFoJRCct+6rMPoxgBnnbS2WEm5c1u4V/a9RZFTPGI5QzxpiVJ
ZlVKqjP7bnnJunOJThcghT13XOCrH8+QFp8GrNyNeQSTycRinh9f4ugrMr1q1w/XMPwlqzxsZCQF
AoGa5ZGQLXRsa1081m8KIwaxEUS+j6E/aSHpej+FOULkir5Hyg5PnokSflY+dEeHIcP3tK4uQpC2
KZCROhdiiLGZ0Jj1azyy4lciM3s2qikVP0Nw9z2QHw8fO4zFjZBeQFr/2bCq2pSa1y4y/2KHBbmO
ig2xqSPImpHprJNAZqa6rWvzLBgbbug++HpR+zyYfgD2/OkXeVGAN1YctmMQflsDmgOvp+8eg8Wu
lQq6FsYgwCc7W5zHKlR2XvhlQHVSYF7JC3gi6eInJIQptLXnyktYZnxCOCVToVyDSz/SWoV7MNTa
l+NxRjDJBC67t0aftVzm0t/Qy4YFq8Fi73dEveyTr5qXkF/93lTEqXE7E6XXqVzqMd8j799+Iglf
yKfRiAM43Vns+GO8OXZhcZnkT/b7twq1WufZK3mIoBpsaLCMzW4lK53hmV/k49WArxDFk5iF16Tp
tp6OmR3rznKT4aiKZMQ6flN2EIgGPjBbvSzKaflRcf+Ha8+HbtuIBI5Nf2D3SO2FSeDNUuSPboWz
k8y51eKd+RKHzfJBuc4LS0mmwrmivQUVxI3XNijaeiA6Ac18389w4frd4ldK/4FmVOVvOLsQ1P7R
rafMTWESfioziRKIl4Tk331NI5gA3R0Z/W8DbVV2LV3gbQYul9Sc63F22l58MbqDGuSy7VdLDOR0
fgrR4eGlyLvLUf9U1/QaSCiWruoGyf5iM3fBnsHVKrBpDFqHQ8IujxtzU5CYVugw8B1CO74k/vmB
YEA2MbmoPh83bf4XYLiJTbDeCe6N+Y99NUH9l1qYWtWwow3C0wnhZmUDpiMw0Or7XIKexnm2MWhi
iL0PSMjoKL7wvLU4cZC/K+ADOFxzolpKybc+7pduxQdgF30pYnvDEPEO6yMFHlXhj4OrVgKjgYuC
yho2HoernPV9nVQhPb2Ej/Bdw5fzXWLCv3TXaxOO1IT7gMBNacBTodOSiWYUjb0BxjJjPSbeIQrc
Ha2x8wpAQuNEBnQ+jD6qApZNLqnIKS9IZXomVHLfQG8XIncmN0RiVoL+YZjC2UQr2SZuUtif3aMO
H8J+z6mwS3f4VYK153WGFAGDj5Qm+/PaWQK0OlneuRbCVtWzTinsjRlXTJr3K1UZVDdxPZ0415sK
WvWsfseIP2cfsNQ4aGXyikGhKe6Ib/PLGKsxD0S2Vx7Cpo2ZyU9H6muT8Yt91Ej+5Dd+keHI2Dqt
VwXxY90PxQCC+SKFQ/wNTIT0ZGuXW5HWCy4c/nhF4vCDtPteE3oYazZjsyE/qi/CTFhym6ExLZmi
9JAZsxEblhavqKkPWh4EybG6Mc6w3n6skims6K7NRSc2jkxTLxqVMifm9nWLdb7QsTtmJug+Wf9e
nWQpgcI1zNwcSOtv82/MKXV1GHzKF0gOC+Vemy85Yl3NIl84iv/wtJtmbbjCh+owl2pnGUXyM+d5
g+XwSgUwdzjlDlZ2mTGeOpt1yUfG/s6UKKV6vOoNC70zNRmGFFXohLfHTsaYX7mGyD7eKYgdqcNH
lCPuA8q0ifSReFF9sVCXqJ+gupxHzS4NcwFCCEZH/ExKmfYQR3PjnVLSq0XWA1fAfwb5YZquGc2b
mPrcjw90X2vb5EZtgtuGsABYLTXj6JWI/VScbD2HoLn+hNG/Bkp/BuiRRBgYMz5MCf9oJppg/MH0
hmHCt0J8TW05UHqrkmutB4GCKNfsURkGkjWJ6hpRCvGOAYsFaGBgCH3oVxua4Q2s/DqGxtFt+GDl
0K68usXe69N0MW8/cRJjKm2TD4a7NIUudX63NOYgGdeSCWzDHcYEdXZg3mvRdUoic3JHkqX0dbq1
FQPk2Vp/ONYsPmEiiNJCCCz2cUxbLE2h04CVA1/fS793Bw2B/X+5pGuSax4xk1bo8Bs/JwGGGGLu
4CNo7k0yGhIPzMqvOEeAFI781G1deHOWB7xbG0LAi6NFjVrj2DrWj0TIrLScbDMkjjgIvn5hG70v
DtLJ3vt5S4IhD7zrUZLaoQ1Sgf97VoF66CsC2pOtloMUr+ThgSzn512SUWmdkeaVqHu+FH66B7CM
/jAS6NLb87J7I8mpORq8niqwdsf7uTL+ylhB312BTZE/8rtnt39Wsn97oZUMK7QebdBotTatxV9f
S2C0tPKmX018q8/9XIz2KF3Lrrh2lZQcsQ+hPM0AgYQ3VS143ayf9FoaWLSX7b2Qau+gtVigUWuo
QgnlxxJrC503bsWmZXy4sDe8NMrmLDr7OL3DMSStTcRbAJkT7PuJWQv5wqnB93IKtoNo9CkJ0nZq
7ZIDgHg/kkJgmVSknionqJXNJRo8j1Y3ArsYg+WPgx1byMLseBvi9lxEFa1P+oY8P1LOeYq3G+DS
cPXayes2cdhP1SddEaB3CUq2UeLnrXiHyzmm5n4d4LM7zUECPg8myRUwIrlabFc/YP2xz3dNQqyx
Woi3LhP9JUGXNxtAWcZYePYWjCjjE+Xqp2t6MQ1zOEwaRuNZJPkPADqMocLE8F5swVnoehPpy6qw
o7bBGJvhYkTlvwmWjFJGmGjflPIbS9+dglx9tmQP3TSa7842RMIHUJ9w4Oy8pBiiknkukSPfVENO
5ujDOOqymQYb73sS6YcuJC3K5fPvURiA80COqxkZp013wN+fKwmRgqybi1ZhWxS/EcxzwZZPsIuN
tffG660B0RH5H3mH391mvTbn2cMtp56icP6r9U8/4OWaSt6DyGwKwXum71t378LNm4RkaA1g5cso
JjIE2f/t2oOOev9/YNvFlKnD6uTg95J0lWgFzWs21PiRd0Ln2jiE1x5eUVNMy2irZ3o4ek2tuY/W
BFiVw8wlAVYc1ftl2E0qgJurmhPiDUoJwUUHOz2L8piF86YqvxmCaxHvaFBiIiVYKlu1JcRY9ZPa
ZwnYzRaFlfSc2lxLzXTNKCLwvWRw0yHOtCyF2245cLW3zJpJO4fQNoBI/tnw+mCQTpLeA8W2/89Z
gJsZO6atriDwfeESjGhmSXX/DNSuY3+3/iCOdpyciv+ES+BeiOsCPCp9x3z4gBUDF5wqwArS57xq
S+oVncawslksSwzg0AA9Ly+KBxy4h/9KSnY0J+0d3RzOgJ1PCv9S8ACWWt2gJxZ31ghINRd+lvoA
DbVFPMayyimjPybYuSsfVG6ejafO13vE1XJ5Ef1RUz1Ydu41sAYB4ja4/E7ORDuuBrRRdnLPmKQQ
TZcOZBRYLjEZyDYenCBer150hV74UHUzcR2R4D9NxW6naiYdYbY4svxFB/lC77G0PmjSppqL+oL4
j6Ts7O5UPSqbBanRN3fz6eUX9ocsXoD3FD3YeuU54eHp9RxoUvAY31QuJSvsTNmoTvR7c1XLrIfA
p6WwMPVITBHDtnfpfvLJ2JPKDbDzBxhsHdZo+GBtOL/4cbwIjjuGrvB3Pi03XUuRhlS4f/K3EbSA
jno75UzQTPM2PNCiXZdMEnwAKe1lhBtCPcVkAueLZrTfCy7KzeRc/2tNeVGdIbaS4EEf2gIhkG0v
W4WUCTxPV9fSrqXY+GixnG9aozPGdBw3ZpEM+7Gy6p/DOWs/pnFVxvAQqiZIePdz1XvXX8R+xvhX
Eeo88sXcXNOE0sTLsu7IFBTphUZiSSF2NkZwyioY/sN2F82Kd9j7mhb08DWrzPRtnRJQfedGq58E
meYEDYrMXi1abAVFgPz+kUhSht/svSlEawDEiEc5mbmHmWbfXAFNI2JXDlJS+gTKU4FK35vzchBA
mHOaatjmM2fQRwOCNyJnAelvel76IurW8VfFgze2vd47xT7WUSgo4uOa3XOIu2SwRdHz4Jw5BRSj
lFxerKHNgJdAZMcIn2byebKIr0dwPx6iF3wC0Qo2fte6UxokvrPeYVTAcP0dFnZiM2xzoldIjFdd
Te9lvgIHa7HUfWqnpH4KfRWWnCA82Izx/lpyCzs8H6aF6VjF1aVmk/Rhx24bKqv4M10Zr04iuQrW
y4FpzNcqDdUQ4rlMq7+Wtt9DLeF0nMQxWGmgCripuJKGWQCMmu3uNrtWjn/ltVQIrhR04Dd1OX/G
J9oVTG2jVZjSRRtTHzCen3XnzyRKTJOzNo6Jw5gpNA0P0ZIuRFx0S4+DxAqiRwzg3GUuU9JwbQMB
mwwiuOPJUG4/BScrwiC/UbS5y+/MU3wl7Ekyjo2hJBTMMFhgAHwSDmAFilM9r4/Q2Dm2hztWhH7G
FR/T7FqF3F0SNRKPD9etiWs6baFSWG6hW0E8DMzU9FkHCNNWdG01B8xbwkfEmOCALvaWYjgQ6IA1
C8c4/NtOIZn8cN3SkN7lDrGgcGfuot9w3+UDv/JJw3pwk1MCyOrM3kaL95fSzk1kwtUyHih8fFN0
bMzgT1gu1BnXTBIH9pORjaU7BffNGMSNeKvDE/gAoddEqcq7IGH5/aK8Xp5UYI21fh4U7HpdB6nF
haLBhXxc3Es2GOXiL8M6w9eDwmgzvTlYBfUPyPFtjQ7bV5v8YmCADMxDBccgNfoSdSGmd6DCJp0V
0bnOo5ABDecUPOiVX0LPdebxH4+N27OOjDV8wDR20i8X5XIUmVA1aZhbaGtradgGTtGrUsBx8ezU
UEcUzWFuZT+TrzrFhs6wnGZlmUWNONk1AZht8IIGWRn2kxaFNDo6ntYxWrkLTchZIIvG0JoUgBkw
SuIHGjQW5TEObLtzG83vXWwg5DW9SErTi2+9g3JQKewLTUl0l+RFIC+H8wj1gB3BO+LoAI7/yzTH
5uth7xGCvyQlF7NTayIgrTn8c4aGTxi1uHvklnkDsj60zjEozRM0BfLFF2tKFmgW/YZlAthq4mi7
y24V+N38BOTVvyuUf5p1dVoSja7LonqVn6FPxyvIOEYsd+ZcpDx2OhnVmdUP8DDQjhQdhB67di0o
p7jHqpaJQFUlsUO0ozc9Zv4nXMVULcwS8Xgh5qovmWKtWofITzSMdjT7DBbKrg2L8UzKdyH2lvqA
/Un+P9baRStM52QXsO3CH7eVtAIL7MSnx3AH93zB8g8wg42eMn7kaM1mFUffg2d5u9o7nx1svRQv
mOVTpvv8NZOhHSm/hJdzOre+2pHwhR+nCbZfzwIkoGeXl+ldOUM05S1Yo7IdoL2HgUn/okutfJIj
Uzbo1Ztp819cAV80GP+S2DtXxp6DbLANZqxZBoRMmJQn0doqCWaFRwpPOXbgIbAvxnteJH3pvXP2
Xo+fiUTgj8bCzWSlUItsusjx2ttZ05wAKlw+Xc9IAuOlqNUb8maGu8D9aZXkby8qfw5bEbGarjyG
V1LSEDqRgcFXOpVsxkJ90trbK6thepnmRwDAk3htUpceawJbWTjfu8jf+QHmDxw+bB+wxEI1cgTY
U6+mBwl/wkU7aYpP7DmX9y7Ylv2OgGAHs2FlGF+E2bzL5SKkTIg5tiW1qpIyGW840oUc3lErxzHx
2arTf6uaEJ90pbcElHN7EIB5ysJat61qm/Kg91/hl5LQbmXm0cKRWzcEfLNbshDMH9vOYko+A8Gu
2G0rckGxmbla747DDypBDKi5x62mWIJL2Ou486nTqwzAke3bL/T+qKonXnLMqK3yk0c0bPzqFSI7
d81WADDcgucKt6M69GX6IFRiy/uLj5gJyB89X8oj3Wwt5TZGW5OVrPkZkCOu5jnIRaizq0aGy8nn
O9j///7yxVBQSUUruvfWPLETtgu8T1DuCTJc5TSELYAGwAqFuBlx5V5+d2Z1W6o6D6365FJWB4KD
NEjO1ioSE4+kZKeLxSmL5MHHCkdqJyGG0cuPemgiTDikJ6gv3Uuc9+W0476bLYeNSg+TtXaR3RaE
41BFUurT5MGd4qZQZZwZaSACr1VhE/kEWqbTeG0hG7asii5Fpg6Q2eftwzaRmCWICVkWRIbjhiuv
X5J1P3PagvBUgnMtRuBgtIdiW3Y8w3PEybgHKSWSrVsPPHkWpADFRTZRt0wGPfCL51bUGe8+HQP9
kFm0tF/phdX/t8tBWcB67u69QUrUhcZHxxpXAz7lTmdQJfUEm1nirKyW1LWPMTgf1zskd+fFF+tP
XNvUV+uZRX8ypLnwIWVotxrq2yHTZWOOKx4ccVcGgKpSTZvotIQxLy32xV+WEtb8RiHYHCiyLTiG
vX1Y5fGeynAPheEpe6JC380NIgPvepF/PkgSLY+4Ar++8Q7gOTAYH6af82rmgjQxC0ZlMavW1IZE
eqn52KkX3B+K4uHOo+0+f8FDSEvUem0lUA2uMwWDsXf4e/zfLodd6otEFfDZgmQZpduYTeBhZv0s
EHzC6QC6s8Y99CPFS/J0qzeJRXkUOlWA0mBlwPD+u6s6c3nt9UTASw9/ybBU6jXOQm2G1TbNkZ7r
BsqRj6t8anxlo1yq3EDb0wVz14aIK4bzfg+PsMWODmKyYwqaLfJMo3YmW16j5ZoCqGxKvKoVS39E
IcFGFC3JPY7pHVzczkmJJNfF6fKjRiFQywsqnxKSPWGrMawDlW+1wBmAROlm3TuBULgWh+0S1VXk
gMtYLlOzpcqHlSukUyyyrb+qVJp4Q9+1ZcknB19vg+oNe8IzP0z/utcSs7N7QbsVqMy3KkmSh/T+
X9ZB8fLvPk921T2P6OfOr6Pans7nAcoMmZTcMNP1prYPVqqBhyqCam7P6YON5sdurKMLsHV9cJvN
ktyKEyHNOKyODCZD9JkpjhLElMnl+zYm9sVNuh4Nqmwa0NKA7ENrRClvvfb2pMFUHSEtT/LxifML
yB7YOvdT71mHq2fkiXRpGxPEQYaQg+KJfRykOABqQFEwD727uFyAMRYhZTYrvvUasl0B0QAIwAxE
ZsT+xJ2YdPouSznkHLAM+3ueqPAC77YGbpIHl7shtGj8CAx2z3+dYAEI+0uRf3KxV3ktqnZJ45uO
JCvzwFvxj9GxO6cj2jRyeWX30a8UPdlix06fA8Iy5R+8uhUDq+o5Z73563oIKul6D86qfEwU39XL
i/MgMw4kXO9ZHftcqVxncDi7atS1Ty9oM3tFdyS+9DNyHUDwGsfYndAr929E1KVoFl+1QJNizMpp
3obegcW9U4Z+xpTmBUXfKOgPLjyouuriTL5rRUrJsBNi6MLHpRDWCVqt6AAWF8iI688Glr8yZiFJ
9itVTbeS25dncummSAqFQvivim6QbEi9Hb0w1khh16aXaxMMHXyxPU96AIo6ph6+SKcALs09kQtn
zylUk5EDiQfOH8CuSSCPf3o78BP9i1yjmtSmcx/44d12GNO8Ar93t8lQzBio9jGZLKAyU05kBLMZ
KboZcktlZg+BPv/xXR0EniDXfB7dJ4CvHd0OBCON1WxhBgXnDcVPVGL4H3yR4Ue8V3zZ+ajrSTPq
8469euLkxPDyrLofcnuerpR7A+JoM7JbuRyJL6VMN03Stt0QpOBE3b0MSitX0VXUC4Is3ga4UOUs
EItKDYMpP57R4/CdZcQUDYHcW3rUikblK1hte2or71VjkmuP95BUfol7FDnbxS2uDgKvE8e1MLFJ
M4egO4I7XIvfj5JRMilOatKDcoaEDGZobOFLSJN3CBqS7mJGlfCXpEXnVcgMmpG1J6Q37uwwZ963
8bGm1XFMZOlQqlNqoWiVSl+7U+FnDGmYTnUoQfrnl4MbCqe9bYS3BYDYOrr84LvD9sWIQGCn6tB9
uL+l0PMjb7Nz9aKqqXOZKni9+quhNVcRnicqaRweAkB6FCfv4xgLQM0g6kYYiaQsw0/wClj7caOy
zjj5FRQu1R3+lECh/kVwLEc/25gJ55DwlNYILj6rOCn3EJXBQkP+yxtzOE/UAfT6aMEKJLr/Gnie
ItflwHUQjRnM50meIchkrk0uc62YBmcXJgsPMvpcbiC/P0V1ZCeR/jDi3DpwPClKC1ldLCTJTmTy
UhKuZHSB4cFpl3MFuymAzu4And+0njcNFRIhxrC9xa/bk+1BGnbvWtBHAMeH6ljyqTGWjvsP02dz
kQjEv2/VdOif2+7ZTRfRqZCdhAUS+lAd+/X6UceozMj+Pb+9PwgCy+P/3a+T3Rp7EXWOZFkn1vZU
M4H1DduqbGtTtkh3YtkYdSy55aQr85Wgd6z8Xh2pEK8ukfpYE5LhZumNJReEd8kyqVgjCS+0FMJe
AjtbFTFU0OlMtjkDvwe+30pSGgZ+5p3HrvA8I+Trn/mWSnJ1JVwDAY+h7uke2GEYYa+uy5k+dIgm
ZzrN+v1r4pf/itvtwOmDaIwFmzysqMCZjjheeWsm0hsszjMtqWbZ2RXmC2Spz08X4cjKDMBltcZ2
bTPe57YRjq+Nd3tX/W9eWkb5K8z7JuLIOmg7pmfJjlZy2zoh2eMWI44rHsGs41x7q3msjokEMr5b
+vRif+KiNPAxuVY2LzreFs/yh1aV1GlmOY9nHeaHNVAtE7SpTma4leKW7iC8dAe4wy3Wzlw8BcOI
FHgMrkgi49n7/BjnbmoBXFOYirwtuN6NsIxOAzwJLH7gUY637K1Tm3gvXRcsDzF1U1/LMegqFoRz
MubGoTLNlA/P8hZ3F8o3TN64M1LiX6u8BQF6B9Q7DRtgN+ECd/Sq/JxsUO74McfaxpLn8SOIZT0G
iDuH1928RKpvZH4eIhtjNeb2uE7tHl/fTFw261lDmnlhAr45v0gZrlj2kJ0piRx3GK9nlHhPaePq
zgOdO3w5nlglvcIRfHz4yLohLNkTJfbjawLPgVcX2RjNbTeN0ThpNeAEPXfdRnpYK0rzEHVOaVh0
OdG5U/mmmL2/pjVa4XZCDFu7/8sSVX5KC/Z/KW0DGnI1Pri/8r2zVSwfyBec2PhhxbQc7wLBpn1n
hL40nuUzsV7icJc4tBkqTpogVPgsZ6IIAffYT12qtNu15CsFrQCfwZoyYhcIjsH5hPxr2UM2AWN8
o8s/EJpVjVTfX1ZtB0p7jYv2Eugz8t0Rj89pxBeNd/itpTOa+OugyCaENR3tF87G3sQphD/Nb6Zg
XF+/fsWf7iiNhtBdCWLnlr+VJTN+0qkFp0udwyAmNMVNnBjJfIlXEnQNcKqHTK2af4feVExmE0Rc
3Mr/I9NdlkaVIJpyANnfwltQcgbii0Zetrq4ZgQodu+yHVBlsW88LuN7R07ogLMO8Pmu9IsND8Q8
pTOYiMFHCpfGv7TwQgT/MXVrewAIj3SgHZmKOhmUiyBZKSbBkVLG5VVCf+djKIIS9i6fE+zPK6uz
zpTkCBE3zUtz+j2ktA2jNcXy/161ct4s0On+dHJHuP5pBfzb1xBX9nbJTlESj3eQjxRbqi0s5fVy
38YhekAElHFDzLGnvpt0b6umUhYexDGm3ZVVFr6EZSMLilwink3vjZfTtO+u3z1mYYSQMjsqlO1R
x9FHXQynrL9yUtnOGvWWrTgkBfckKs7euU7d85CHzhpPC9v3jV6y8dJ8Kc3QuMzTCymcv5y+nAMf
koDChLx/kEwQthd6BHGwPfRsxyDfmeMLf8qmE6n06a37NJbkEpyOEvdGhOBvwT6HXtU9OCmBazCY
99yvlH5kvnzxt8jmw7D/hFlUxySuwtyWvaOg4HOdjBR+zcJKRoddc2+4a+DVrTBD2wbLWnJFl0h/
bnmbDIsXxbAxfrR76HPZiVrI/jfT+09oG5B9P1k+/wKJv4/NvRdiclSDOFa9yNlHVrranZaWSapY
M9Rh6rKeeDjh33MF+P/Ibna0TWYJAlUSggijgyyURw57jFsbVq7dBauYn7cUbzUWmMb7umIL2Rfh
SQohDCEeVMzfltWKG2NhUY+/8p6NeosswMsd7pe0XBV2j4yhh4NtbeqGwahIltpFDOvtdy50aoHt
z4v+sn1IcncROOAm35yaPvIZvRLi9BL0OS1euSscaPJMldUDJ2NDoPm9aYjT7TTN61Z/x0xdjXLb
yINlniCLS8CLj6TUEuFBdNTm7NNE2U5mGLEouD0JdTAu0WLCDzJuxFwDzdG+26oftOtReGV7pgbz
0/oBmLeud3ylDiu03dmRgAOdZ5MRxpEjamk+YGtAsPUjrSuxrkZgg9FxfJmNn4QMszyqRe7EG6xE
l2CR3HqtPZBTfb5sHkM2ZNQPtAk7tllfjLnvsv7fvdxR+RoN/28LccBuQ8+VPQA+ipi04aCe/B0M
rwm/wKQojehF4/h8hyjOJhQiql83cMzbCv7r+pXAhZyFISKmiQg0hhnGPgyye9nlHv29ePKE2lKT
ygRy4dykgijSvH8LTDAjTJFlelFLcORgLnaWaT8Lpaauu8Qt6IOgaX+FI85bCiMFC+z6RRcRgxew
uY9DrlumwNWO/0tmrCl/6p1LF4okw4gYCQ4GjoZ9Mxzx6cbAtKoMsu/O6j3RMnW5xaFpdv2iZPZV
MZAUF+IqZy8FmfBndioRCWu4Ce/IxmmUCX92lp0A0FRzDKH2wCTuHaI/D33zkOYuSzSmMjhnTG3d
RbV6ZxUBKMHeBwIDTzeDrmRGfsHR+iUNn64RhKfrzbjyfckGQL5JB+3LQoo5E98LpGVVADVWmUTJ
n5C4O+2N6vN49SN2K9Nb45cVIwm9KQcj3KBNlukWFOECtPUGenqX4u1s1v6vezDybouUJiDsbD/T
Ypo5RpoeP/Tq3qZn19bmgG2HT1cpqWNidxpQpwkEei4xWtM5CFQypuX5G9GwtZ3PBedJVWbHK96A
0mH13dUMYGBHsJgFacWvLy8A9HrTKy6V9yANKy2TuYDR62SarDph8feUKuG9Pmvb06mhEEb967ST
2V9gllxB9OKJ9AJwGQje5mDlpnIXhbr//W8AxJvzGNVtGnYrkqrc/Ia9otpQhnpdZ+W2iwQnOdzD
LD87pt2gAlAk1fkIEd2sZ2F9zSy8zh5qTnZm9g8H682z+4Vg16TF+bFlNtKP++qqJBcPCMU/gsyv
jucZm90lQPenvXUfwpkTUATPcpuSvWyyixlu/fLhlAngHbtWy4Md22ENaNHemoyQvBudEOAA6DYO
xSLe54LZ47UgkFjw1sh99mYkhmrEOY57Fzny4A90mlv8NAtiLb5u2gPTqdoRF7HbMigEh/WFxIdB
nk/m4egXkkYCW+EQQSPBKS047UFir/z0BEcbr3vpYEbAgoOz/e3nGEo9IzpiC/1eTx04JvKwnLSp
795Bg8s1T4RoXnNagizxMtYkROBGG4IQsjCM9N+Bq35kerFUjxhXeNO3sOBgXCw77n6H2Jh1i3ei
Q8N2/UHD4RiuznWbYj5JUy26DyW/AauciJdrkuPyy2M3Ra8nzH1lAraWD1h5TFvIc2oYov23Y9qB
xvD/x/or1CMTxrHqUwvP088njIjtturOJdwJQmkj58jHtN2f1eI80O0j6bcKODg7TznVGLGxK4cz
VSTpZ+jO4JA0uNlDpFreWLp4Ftj9uZUD+2zKDvJG47Is+hw3Zi39llV+NREdgXUS49oNqOSCyZ4T
W3ufVMJ2uNAbrUvVnCg9NBncqzt+4uTklmVPHQNagWiQ68JD9Ml9F+SyDP8WroPj7reBM39QBq3N
Hh1aRIc4vpdwsw6hBlJADSyCnJXGF//xlDr10gnC5+1IFvf195TcQ+pg9xe1EezNwcW6G/0cTRBu
siXvwjfN8rRSYGTIcaWCb9uLhRcqzGmpiWLXXKor0K6yxDLMbvnWAZdEBulA3aR1ed3P2n3mGACu
mBxyGyCFgYIVnpKfp6v6U8EIgSMPvKqlePRgvUndxvJcV3ddClmb7EnwMS/t0CL2Gy0w+r+BaRTw
4JIboOJlUn+AV8C/8f4d1W2VHV8MbB7exSo6/fj3TZpWryFtcX54JUhOPAF6v8T4s5t1zuVoH2GZ
mCsEZ7UVlac8GszdnNauoSNrwFH82p4kj7x1gsLk80M7knZ/W66dzFRMh4rsiI3FcZuHzE3fkl7H
zsXZYcZEAx4TCNzNcIxD+YknyI9+U/94Cs2R/u9dMR/1aEMwaSIdQlSZa2GfhjOp1tRlfVJWDiyS
AMCTloQjyLxJ+ax167Fnce7th8k4dCJxqtueBRZPvzXhiu8oa+Hq29XfDXZ5MxJrbZvbebi5Ockb
ZBDEax5WxkSUueWOB/3hgXtmZxHCQ8FZMfJZfcm0V4GakgN2lKpEK+RY+xJSkB+2NpseJuYR8q2i
BBv4tqfPcwWxryzJ5FI9LNL1JOthp/BuGV/t6PJDBo0Z1EV7HgVd+Ig5liVaaWryCDyG3ZJ9+VuX
79xvoPtPqYKqIMaPSGIIHxMu+bBDL7zCjrw4uBOG7oA+tEn+5XxyoMb/QZadQuXEADHTpFmdfpnc
1DhAKEK0WA8rf5PIlboJ09u2SMLIsvRoKj53WrcYPAN3xo1xNN9w9sJcxWSgx0EeZpXD3QxckrQP
Ekg5p1mdqmqPt6cgjaAzV2do2d1Y7eGPFlHttJGZOHtS6xlDA8ANOsBdVmAvieGxCGoRYXHqpPXf
EVihdTABPuql0sfTZkwZ5iS33SNdA9S11r7EJ/qlxYaFuxs7hYhj8taA1+oHeuybOkX9egVFXzro
4Ut8haPF/x8arwY6OWlnvckcmi3CThs0tMTaFdipii6h/mfvB1VGlXFYPyjcUdvBPgePOAAmgL/9
STVNnzXFbTykzIDKDQoc7e1qMGvgnwJUj1LU5K46mgBQ6Di8XmDc1XOcCFm1iqIIAAIgJGPfUzjR
1JeB9kXX4oqGqrsqHZTf81hXNQYn4nZigW4ZeE867zkUtm1Wc7W8WSv1MY3/c2e/JHlQ59OzOY7w
nz+4mp1AHpHzhOH8meizaT0ShGmqunOJbXSrf+X2Rl2MzTeD4gk2giRPeqys2mU2ZUXXZF5AkHuj
GzXqNfdgSMRGWPSEKR9AmFFbIuCigfIlx8h7a6ONTZnMzQtqwSdwZNsKROaUZP9FS4U4UGKj1gDN
GDpgSauLg4HVq2OsHO1/AtT2iy95rLn1+kzBKRKsA8Hls0Rid2zRvs3ZxStEat/d043OZVFoJU6h
1sKrU3IJrO4jsNpi7+F2aRRjykeblGjs6amR45ceo4sapua9ZhZ/BgASdr+VJeqpeqsOe0jNok3G
An/9VcnX+CKOkiQoSwCvgZmZve+CdjN9J089K+TDanLtpGjJ0GbpN2HHV6JNB3+gk40wCrn50G80
TRzTUhUJ+Dg5x753w5cy3SswJSnhj/lJFpXSmoEkHKXnaANC+W+s5S3cemT9Eldv4reBedxY6L/r
LXIo1jaYbmY5wyCv1Wxkw1MVa1V8oUb29VY1xPmB54tGQ26usycLrhcpTxgZw/g3BThAYSPWutG8
gjLfR7W9U8fpKLZHtc8FAiMbUSVMsa9cKbXFZANymk6E/+qmHJgVGoeNV9lTB7KvK2trTJ99l0Gw
SJ04rMzSurWs4xD24Jcc/PDMGakwxrWh8AqEqivyTVZik6MypnlyV/Q9vPJ2sIEMTTa9+adskyMa
GHINK2OgYfomIa0tnPI6ZOP4WfRGTzl5PI6s14qJKmwQczp8N8A2gGHPqW7pFuWvmWhJmnQp5e8F
VFu88Bam3i+X3oNl+XLGD/AT1Z3X3BgMLUdYU7dPoi0AHztovGw5ps72DOdMnRENghUqB+VbvD1s
2AqL0UWVJY4RWSIc43+vtllCKPd6qb0WynZP+Zb4VOvmE3W1U3G3BeuOtE0g2RyjeIAICIzPRNph
Ks5RWVVAsyQWC4qfnWFcpVDQRXNseFCBH66gdz43MGviD8phf6OnGKIPw5O2QSzVcXpnhTJKea0j
slkBvZpmcqlPkPu4mwjHoqOdJ41LkPcp5ZuTwx/xjR0xSoTXxySRqLqWFpyGfq4omuhltLnKesMW
9P12xdYgRaEXh5UnUfBfqnDJMM3gkfHZQyIUp5qyMJN/sRvEgQjugfBP7Ao1pcKfx66HP4EYiHmF
GWf66VsMxndDyz+clToQPjvqvO9jNFuvlvHPOWYc5Q8fKZ5jYBgCOalYfMglbnl7g20gSe2Ru4JW
EiZ4xlpdCyvw69rYEM2BW9aKjgUNYo+b7KpOTSXqZcAW1CSGSBj/ZnN00AQuPoB3RJdGW3SXyMlg
1qSPjoKWlDeRuxCjvp26V7u0xW1LWLBcp883DqhXHnHECX1zmgz1kF2amJ+10ppHqYNhkRkPlrWy
kDWzyTDGjLq5l+IWJh+VcfuqHeJqgrxLqsmLrhMFjUoNXo5MIFiz4GQ35yrQ4axSr7T0cCtvNHm5
LLNpMWuG7WYdggnBWwY5xXboLbk2PUoBPkW4ux1P8uVNOwj4C0UiA72YHXOOLgBs/thHP96K6Qen
0ICeeBsub2/FEhidQtnb1PS4Li2n+I576b503cboY0JEsDbddcpdSHl+DDexaGETgzibByedd3RX
A2lHB0kTAgYxKcVoZbjnUIxfBycnupOdMCf71Da8iyT8xrsY+edlJH2vYTppH0e/yzmVPkMg3Fbi
dq4lxqBK8NcPLDWC2RswyQwMWJFeuUOygvWzTsb8CqZ+cDYPmC2ht8yalIgkU37gdCGNDzAmiPj4
H9QT+2jlQYh1ZW4pMGHnJEuXbe65vttav6+Mop6C99d32fHZcc6Fw8grfOU/xJvQRzIvXHqnVLCy
VA6ASRp0cRmX4lDcKDxR9ZNGt8g4WZFR77HeW7+/kjsDTe/ttBlVQ+PUDkhSW6L/JEGuZqrKv5YE
rjGLxgh09e5LyOgFP16UKmpRC+aloMg9k8eV9o/+5nUxGHfOuCt71MTgDJ8KqUdHTrSlo7sK6FDv
w/wuUCLklFRVNbLY1mpnVogt1TsX8Gv5hogQsz+G4nKf2L+9CeEPt1lhwwSIOy6TtAqCgXbhKmwt
YAcMqe7ZS5R+5IMqGF8fxk5Hc3tOxjroEE5nPgfJnZftUcYeZ3US5r2HdKejOrOwUwoDmmBJj12g
uiDlqxz8Fhyq3eOgn2F5emli428wfqf0IoYd0v2YtofgDUZZBjaJhGtBzkApPMiLB4TgJQWAQwkk
xz6Ig3aSvl/INVZkgYHXnNR/d6x6DG2NunMkh2N4GpKZTh3cuZFt03lHeqvHMQ632GTVs47psHwg
F+58yQPZSW4lwjCuIuaVkuhvj1b7ezOarDnQwXHmefyPfbdEjsofqj/yhnjx6ayW73Gs5mIKe4uR
pSD2LLCfSvfdsIJGc1+23A7CsmkU37nYqsokTMjjKoOhYodJUZKiHCNRVLNjSGWVcykShkmjJU+5
QVMPCoDAs+GFsKDu0FvaCrWOmhxHVi4I5p/6DEfB/4wJvvai+FvB5KjSxp9RDcvrEjEETlroQlst
oTd67p3ml45f5ReJjabSDaiGgyRrlH15BrLPn79okkkQNreYcMLxQPoUSnYCHrYpp5rABXdunZYS
R+pj0BCUyhXQsNwT2Om6+d2V15Tz+JVtrTxAfrusG1T50/FUZWtH/7Fs9nHhy59xJ5MgfQLrl7hE
jJ+/+jPCzoEogxRb2ayqIAt+0CELgL8Cb0ge3OPKNDqc3HQcc1MjbSCecQujsFEghuFfmilNQpZQ
EsVhyHCCGL4m36YASdi+oh7lI/iKN73tB3HVZj2u0aBAGQkknAmIBZUlkbHKQLG4wF8HEw+SKbFV
WtjX4pAhvl3cxi4OCl0kI1pwv0+louG2FULhV0g4DBuaYBnHiuggCfnxGguWQRQtX8tJnGdgs8a8
iynkoCtpF4B+bHsKam/UVtEFCuLDc/D4fPk/BkbV28gmYFFXMq8UoVdSvhPrtxBWLqQGqPwBe4UD
KsOmh/yTGc91hRCDG0RJVbezRj9JJyFVhSoFuAxhps/FLnt7cTetzvmFTUhKe6FzIR7B7pjNssNN
7YtnaCAijx5686zGT2PPTTrPKPJOkeHnC+uEUPkdI0TnvSvMH9HVTwDVpp1hS6iZ9f8oEFd4KKCX
O8lfUACanpX+QXjOjvZTFixIFXWy0kguONPI47TzXgmtmKG6Sl/L9BaUKDg0YTf6Yjr9z0HUYdNQ
4LsMqKn+mFrnb0wLGHXsAB6imcjT9HnsWXEUXyO4orE+DMxpn9fixYJrg9VLEl9lD2Mn4Ob4mB+j
oDANUQihYJsKG3K2AwHGU3HZYE5E1Hx6jY03jxY9sF+77of+fUvLOn+qAok8KaWWmweT/wyq7zNi
pPlSbnh5vUuOT/h4x+HZoyKrkNTC//TNBRAoIDuL9nJ8CLtu2cz0nsukTUJ2aHm/1IQZJYkMtMHc
z9ZHYrTsNlGzHpgdv0NQPbz4gNnM/i48q7kH8A4EGP7BYiWGYugeGWufAid10Qz22k+cgatYWi0m
ZISlvjeRdVix2uU7pJFfhvw3Xu3i3gzTgAoWaYiMqRm6uA6RzoegbAQOH1NpraozbipDEOaV1V9W
+/cH3V3aGuAeH1QTjnl698UGLHVaivyjdW73BDbaArf76hWzTCDuHShV20urWyniFQX/VKU6wC+9
GJPoIHKRlguJO0LvujcpRdn/vMGsoOrqLgXxClsEaE619FJ6iThT/4sEskVoHnI3JJeZVkNoKjMn
ZxAkzMrB9Mc67QqElsvBHidJvE1fV3HxS++00xl4o0rUpbuKjH+0mF4hpdqPEf+7L/j+75BlJt+M
PXEwgfJeJAYOuNuRy28HjoHtSX4Lly1FAS5ms5KSqhew3cb1z3Au6LEpU8wHEgxkMNkvMcIkXKpJ
16PU99KBnxG313H+UtUaU4Mra+EZ+GRV0TiE4uFwbFesnYQoLCi6T3NeP0Lf6g5OP/3emKEhLkmY
yaqhg3VnIfMbeCOB9Dhcjmlmd/o2as2lI7bZ6aQBf3Jlu8F12ZtSk3Bqeqxf19+zmWcyx+Kvd719
t9uagq35NQRuNBism29g7wxO0s4uCe6FdvTe0h2mjwPjJ/6hhos1srIon3n/cfdn7dKEogr2T3FP
Auxmo+DBlxgYd0XQiUHv7dtRXgdE5Aie1lOP+qnV6VHyEyc1AWRP1DT2gzwlCzup3D2ADjjafby1
06PuKPs0M2sFeKvkCqUmFvf8UnosH6uYy1QbWznIHCrG4A3ta5OdQ+AwbteRvpX9CqRKeQEpyDiV
6Fwmrp40+D5G/T15ap1DTCbVX+A+eNwyG/489f0+EY6TMH81XU8bHRscJ8x25/jGcGifryQk0uQU
CjU0D31kRsE53rQRP8JreYmVl6nE285l7BriglsvvsQqiKOJX+aylXAJlM3VNUEgkr00aDrhrDeT
c7Lpr4lFEMvWYzUy0XfTVlqOyZ0hnPvLxWf51InVGRZLlhFuAovwjnhGo/kREwx3VxAfv6K4z7MI
MZ5Iq1/MABJLt+LCwrV6PV8t4H9voYBk119Uymafwx4cod1pYeop8hiupffd1u1L9PzVWLvHtc4h
10iIwo7f/CD29328r70r/75f4rKLsjcDxOivkvfh62UDVhoqW0ERUbcUR1VPGbxz6/ueiayjYqny
6I13lYj2V+Eg+zO7851Ft4zD64Pv19kgLLPYhMOSxMP7TehGUxQNuODjW3mrgknKw0sWkIRnjWLp
5uHASm2+j/wP4x0bSgxmpsudjmxWLTIrx2CG+jx+LCY2bujhUMykKMMsaovHeRsR+lJFTEwAXfOt
PXWqZ+o+fQHNQ8MT5lu97/VeTI2LBgFB8j76pbL0VifczBBSNoJoXo318b1cs3P7tMEL15v9Usna
DTdNRWR1LkP+h/NAOgOizclyy9Ht6p+P4iT1piiIhgcjKyu0QHT2wE3EUB8MVOsZz71TwhmC8u2W
AfOH5TVKMNzSYS/YzJzDcxzqx9tR9Khhe4+yuu56ZVCAOQzl8S+5iXE2NMXdqo6eknstjKK/3D6h
VPiVo4WSoHVSqcCNChLEvIboEzwhBkBhBywJS6rhN/QotwptdZOh3yM0vmhSG/WxTLbjyVrjp6od
wRibLjpw2oV/a97nOE6VhvpiEwVLtV3RVrLHwi0F8Geow5lRx422z3fi81UvpSW6k6+54fBXKRw9
1TjND+iRiyooqFwm1/28tFPLMpp7AmhCs3ZxOV+5N9nuXG0wiIKpw547cPHRgewitbJQionLhLN/
mw6c9dm3L/b6qwSSuZR+188ZLGckQgFcZm38qscdM8f8lOgHt55P6QwH2hYIYeXbw/kGDnO6seTA
sUDoMTWb0E2dZgWsAIKtpZLvdSDAC1Hnuqny/SWqjRuPo1fnTe8FfjuB7aP8uOGB9Di2te/chUrv
Nc+rNi19qB0f0TRO2wf967fFUoXWz+yUw7F+olit1ipM0SIHgWwdToEeKg1GDCIF3Ga87KQg8v4U
C2oh09BhylK2UWiT+J/k1tkK8HFfXyguo1iOrUJjYFldoFYl2vF/eeXuWVgpx5s10WyCj0h5OOh5
2hzJXj3IyQ7TnaDQOJWbrMplYfvSjBzxH3xLMo6A5mcW9uCzc71fX8Tqq/CzzNX6+QaruxUod0mB
hdFaxMQii7cIt/6IofYr3ukpeXYS2mNOo6AzmUH//3j7FjpqJaAG2T13YYrJIZHAcJgCSYI9Fa2U
dthlVkuvzmUCIt3As7Sj9lJZyQAHFKqJf18yNssE2dyvdSpCShU+gcTjWZQIwoZ0DJyn3TowadF7
fn5bc+kIsLAGjVEx9iy4uL6K2aXSUEIdhlJY7S6q98AFoOivsTSQk+wXwDxWMcNoYbjm1RB6/Sih
oPu8f1PrxGIV9jAZiAgJCw1rkahZjrX4xQNaPy2GcJTqjgGw6zJAwhNpoNNspA8AkUPILGkKRXhc
36Ix2xsCLwNqmzg/x+c2QU/tzE+d2CNOikwPsKZ6D/NnZvjNHeQwlvSaYs5p4MlCgVGhX80c9sC7
hkLrcNmG7L+OTYqhX8f/XDD/ViofBlH8jAAnMS+//1INsRn08JR921hZ9f1/toZQavB/RvTThoU6
EW3Z/2ZVNsSDLQSR088oZ86Z3ducZJnDvwDQvdTKttVCKij0UoKwIpAklcpYb5XQYAikBlWmWlvY
AYmEjOs/7eK6O9GSOgANArsLBn9yRdT2yUeT3CknN+aiR/GqbfZHXYAkobwozh+O9TYuGOMSHUXx
vZ8flhkHwMjg017Wr5QYcbwE/k8WMRtjsECbNFeSqq/FI4pofb2824UdfFsqqrpJ4D8b3FQgZhUN
iCM7h+Zq5cNKslhqrSTmaoV2QKQD5yUKrS3NMCADcE+Jgs2nSFI9iafFGuq8bpJtLG0G9NFTdWWC
7qFTq4VVHf7HmIhjAjAhknzhbrl9HvW3lbmBTL2nXh6k0wSisLeaLm+YE7mz3hSaAsDC5+7QuRh7
k3UmUWkCDzzpI85NQIDrGtfNdHAQUzB+aemGSUiCriUQaR/7xK+Pq6CGYXeiLNwIFKunEVcVsoCs
jAc3ErZ1ZhVV/Q0jte+n4gLbioKV8Eo5ccu8cgSRYOXcWQsLMDhNgjNk5zszr0v2pUd609Yt+/d3
an2yh3hDcpGat3OD4rOoWVWVJdw6hNg3ylraF4oWBTCujn4OCH58skX00z7L9U13FDBLOz6NCsCn
zryWfQSADZxCjucf9fu7jGwDMVl3Pk/Eu/E1tkLHQlY3cA1qyRmW1degd0qh9hfzdnyomx2HGzwF
+sURW5rBpkWwA3+XF8m45d/MKYb+SiXcTVIAq/mRK5fdSJwuDUL6kqwxGNQNqyhY1o0lhSdCA3cQ
Eq1ytHrFIdz8+YwwhwVDLE8bYhtH6FV/e4otkKEHZ97b9B0RRlaiiAfG0nYK+qhqm9TEVSI7glls
3Oo/Gr9XYrCkiYJCiuqS0B+sqmzuh09bQdMVVB/LUQj8oqvYFJkGRWJiP9UBDE60YASTvagTtEyG
6P2T8R23RxawRV4C8yyKvyoxGS/7fZAIbGddeDLixFXMkfLrvr23MDEiA0racYEfKWWAUdZbQcdG
aVqFnbBpA0E+sRAnCllWOBGDHM2ggEr1u3uCeQ8qlHKkeh6kqGoUZRdYXOmwBfkj7DoclxCkQiX6
CglJMKQE1L+M8vp0CqEIIWt8LrG1CwgXIB5CqWpXNlGeks+Zy2Jrx7JygpCx1ZtOz9Imbg01i7xi
od8eHPI4Lcjywx7Vb48KDoGwjIQpkUo1qIBIm+OT5QlxsRzog5pK6Hqx4HLG1xM16CTdi6QbLg2m
wrPetw71sAHzZiUl2NLSMv//4YTDPOZO6Yo2PwAJGJaaM3bRKmpCr6mD9WkTypxejf/J6l476y7a
kVFMNAQsbqV5mkYeXy1qrzz8lU1aU/61v5l0Ap/b7W8zJAcgN29mTpaFzYdGuDyh/bakForn6tNX
5BvJpmVV9glAFgkcS2Nr4tXouP1BXAmyAGCd0pOp9oZxuxapii+HxXVLK6NH2jms6UKoEV5uBM+o
zczv6+7bGPYISGVFq5Pz5+IiX2RKphfgS9NLbl0io7kVXzdFUh8Dgsfd3pzT0bQ3Fb+kn0XYE7Px
dkw2SRyCFG78orp26dET0OqwiAyLlQx1q9ouqn5hGoAl1F19r/1TBK5DrXNLXFHEbj3Vls7ALcCO
aCWvu5mNMxT5MCpJjruVgq2MDO57TSkPx69XDOhxPPvU+xyV7ZhgYjoEhg8JMYN7v5lL5eT7gQ+2
mtNISIT6wPjiUDtJASFE7OAeBnMvpxUZzzBgqnpDeJp3G1ZcbQtQKzq3XBQKfqSKcfSZEXzm86oG
JIcdmIvKxlmTFa45dF59DLQ5nfxaN9CiFfz6fxg/sjc7JQw5hLmsjjOafer/UbFkiKKZOCX6clCO
S4ae8pvZOM1SyPDauMtaVyt/+u++rU9Gss0jTow1Cd3xoQ5hdThTclS8VKlj6KX6W0gcswoKEk+Z
D7+isPG3A/6LJkZ7IaxLpUeNWEoLl38r+Jb5O0X3edbu+36BKOhZn64LGEZ2glppOkHpid+TXtK5
mZzhTvzAOsJ7v54LOjpqU1MhkZTSktjvt++XAvwdg7VMoSsOWSkURyJkqYp77DfldkJjaG8JyFJl
BgiOcL4ZxAfiy2Z3+YnpvqHBOEsLrpMHPlJmUrHHihOYcqOICl+Aw1dAesgXsxzI5zu/96LJbEow
u2YJUWDvywOxu6AfadBN/UPW9WuJu/i3RKYRpz0H5Bo9tv0xe3DrULtuzZ1u/HEXz5eLbRF1ItBM
OfWHl7y7kaDLgqePcH5Xn/8uzcVIUDGOfGKbfSH/ZIVC2NO5Fa5PkB2k26oEEyKRe7qpuXARHLhy
q5NVbDxaS1Ov4BbYMOxomJvPnOKedqeIM8AB+ZT0ryuypBwgjuV8d8mHFWBzG6gJFSHCaCn0uv0p
ASBPHHN8YntkFdm0XFmDI94woZAtzO8igIEAv3T5GV/NBfMw5zSaThtQ1AVxpUlgMsM9KHKBt6si
nXnixmIjYIamKYNzcwpdhVE5InV5IgkOp6ywuWNkQ7bBBvoQcoIlz+fcP7QjOBhtILwUzQRQPmrd
zQzX+3oVTmcBafudlsav4ZvpDCABOxXV5NoGg6aOOMMN0G0nHo5402I2vdsC1p4Qno5C39ONcXIX
rUsDJm47l2Z5HrVh5XY62LtrEcXDm+5unnSYZeOji94oocgMYEkxHNZok+HKt5OAhLf4N0GiXIyi
R2OgMiPxXvnsq5V7DNo81pQECP2b5XECzLf8xAUy2o+g3fV4/CBfbEiPWQDxXl19atFRL6oajY7p
K3+XUr4g/YG8+ogbYxXUVwKqHbXONkJeW6yrJ7EkbPBYTOE7TSuSZeRrAPE/VjJWutAFVH+7jnU3
kWqc5beurpAc8Q1BeOvG+18qHmgQJEz/T1KIFK7i4IidF291gDSaEkOJWbqcY7/l8B9yoxuUX/iU
JAZ/nUdyDIwY6xZTt6xsHlE2ByZ+e5SGLAjgwEup8XWBjf4eO5WcC6SXXKTlmlg6+u/xcSi4t93M
/tNrVbZ03F2tIRMoY81wTYYiOOspQHk4GgZtuIMnX+7yLQmB2B0tGXuaYu8+Wmc9EuVxWBZF0ZtN
4AEkICuAWI0hIEOtGYTswTNFzfDqbrRSpbZEIPp81lq6Y0k7T3FZv02mygkCQ5meZOtR+jiHFf1N
IYj95Db4oZBFTcLMmp4wGpSz9IjmUhS+S6F2P6wHVV6RWRqz5yKhTkv3XnAQk+iiUuZVTuLOYjwv
MUTpmVGYxSsoMdoyH31LzxLBEmdQJJM9pTrS43cCkg98q2SNK/1xLiFqz8xOEiMgoALNVZrVjftL
YF3Xk/S2X3KqN3V7eg8/NrGVhe3AV2Bfw5aWSahXq6CFvPxMdq/MA4vjRkzsupHmngRjigs8ro9u
0WvRahy1RItU3GWezxZu0gRok+ZXyBSJVsZfbnS7Vg65CuJqsgVGjr/4lKtBjBWYkEAoUbUyHBxy
aS8mr3QTT2rEwB+8MrOWH4YhBlI+mK3crqG47GQpgjFrkxs7eXMnlEBSMeP27oGWF/LYkkuQO2ee
SzEDgaUGvps/i27DN1vfuIxZAWP1yfHEPkuJdHh5zTuNfjQX5BINvjrHR9/cvoXveIvzgV1RXC1M
uLx81nJnlnDGxPWV5VsQyduf20PIz6dxHI8NAq9rG/TiW3rFeYIeOvwzqlY+Wv3yXWEkFzZAWClR
3B48X9n01chLFPg9Zgi3R5dThRocgdpWN3U5iuLU96QwOSpT2endH8704dnoGr8zyydOo/MubqXA
M81Uz+uv8Em2kWl6DQ3VTadzajC8LPvWMIV63jNgc8cNvoyCdZwM3MzlzeSB1wVTsbiJskeuIYMj
BqG7UEowZYxov9ep4enWDIoFH57EmGXd4Z/Q9QMfZbrWkGtJg7XCEs2oRKOLlet4fOclNwC7cSCz
ShfeZn20LLDZQO+eqZoc4lPmdRh3Y2qkLRonFVGbX6H2jRdLlVm+JIkNa32ZDNtufDij+OvCCjzY
dK8sV/9iXZCpaH1GMwuYYeby9VspxH5OK4f7J2Ea52Yy++3CXxQ+37NhLv45m+mZzLnLriN/+p5N
qknginiZVl2vtxOJIQfR16Fu1Fn9c7xLthtuejUgQr1p5CAPYMboq3n/r49vXwvJ5aqN8I2n74XP
aYap/eFBrtl5gOuqiA2q7u47s3ZRKZlkcGb9VHQosdC15XpDBnIG+8AF1HI+YC+UVPOQEIniJTCA
B334jG8DQCnvWmXj61ociXBsNEvmWeeUYGis1Pw/nOzI8Aulve0OdJKZ58iplDczYNF9fe2d/wh9
01kbRhyY2YnaG3Smu8oTx9T3COXd6FcqPskvgzvLInHFMvdJ+dHLhlms8FGl8ah9+V8vUb4WYPa+
VFQUSqTzcYjddK4wKfeUbp6ZaW0pygnBVzZqSCWyAVVJMX/Fs1Fn7H1jCf4TWfM2UAYSe7xi7QQW
0qRuPqf4Vpw1pgDMkuZLcw3d1dZVt4lfC/ZL54K6cWZhxLuozu+QUSa7aPkP8YARhvfUzvhc/7Qv
lRbfMRq/3AThpCD7cjG2cwHjSafdCtYfELmZA1TUhdZsOyGnpJ3kL0irpUzvhw4knwBkzXnPTUfa
pACFTypPQQfgN91YpH3Py6kpOVYipwuC7ydHTd17wzwrancv7uSvfU3kdDIYmog1ARCVjKACBteZ
vJnEAOzFJ5Yvlu2JBuT8Mj29s5Umcecns2tTvacY3h2HK0swt+0AqsbF1BXcEfhz8UWqdRMIFLjE
+Q8pGJD2adzQ9LPhbu6v1HeJGl44T6N93X4uaGj+2dg0B/MxIbYoB3+SlqWOlXCafyBXzR8eBBCc
HUIEkeTZTi9xP7uvpS743gXADDJPL2Vie7THZDBsWRyyo4ZjCHvHe9/G6Vz9Okq9bQvO5yJoe4zG
jFFLS3hsk2ndruZA823RlwDSTB4tf7rKvf3KJHqd64nFXbA+bqSfAOersE/pT9ewETcF99WuIAbL
Hck72sgUlMTfFr5PxFGu2E0a4BPR4g9r+xiNo5zVX0PcvMKOpyt0Wjit2BB/Bs9jyrxFr7ZQ3oXp
Cm75rXmCgv/F9nvAz/9CL2HNwaBj9J3qC1tpkgIbzMkK+eqEGkf9b+WcohcgSc2omtbC3XAWae1r
qDTRChpHMPlz2D+i91AnPDMk0CHuVK8Splan9UeYfGpQR1xAsGYuBgQKpAyTV8AsJjsvVHDDGdAO
Gb+FR6CHXMaJNsPPPN2cHbjg+SXxBbS/b1siaw2bVjlJeNpdknruoihbIfSo/d7edIGb2NJIoeXb
Z3GLqMyV/6UlZliWq8PdgudI3uXqEHs6Dh3e6Iesf1OWZ2s+XbIRBBaP1iQkRgXzVevVZ16iY8oB
LTMYtZjpjmLiIdp0C4C0iqeCw9mN3+pV231qp9f6uqgm7myaVd4PxT9UU+zAZkCbxNd1sO5uA/B9
AQYn2B+Xay+SNQBokKH16zpbGGmxZz4s0PCmJdOtb3G8WfalfIwCQ8fZ/hFP9LkJH2z8s6HUjR+V
mijAmyyqTX/wz+pJYpjO4YxWv6ZOl5d7j2PldHemp/kX/aVBCSC+BmOYe7tjdLd7CST9k+UeU3rJ
zClUV5Oqou+mJskYSOAyKiyH4uX/E2Iy9wTPhBa2xtyrO+MNkdX8QZOeNDrP+RK6hLXlT1XhOJIq
f+K8zlS5tFwNssjuhEGJ7L+HIJaPE9lL4ONB20Bj5rJq/MUFsdAemNdMKJK8NP5/F/kLv64WViN5
vy4I9RvbbqhPgTWecDo2kO3Zf4MPYKOjh/srbj9AioD3636M6qPrWweEuuCJvT2MqkT6KJXTvR0l
/fL/vvf3Z1dr0IE9CoXrneIJxV3ZyxoRMpF1D0ykZ3hcdCwNJmRGmOJFH4Mr/BRaACkwbHaYEyiu
cQEl+8gtJM/v6SIAeNu1dtdYszUW9QAwyRSHFEvwQl/5RwuUppTm3+hAb6PeYvLSd8b7SKAW/DLv
JmDatYxR9IzCOfnmX2qVFdIiO+abWdDF6Px8qtCZwfYPDvARvI4+eKJV39l6NpZbJTN7DUSLN4WW
VFZFkKJjQo5wEgBW+ZlvJgbpJj4Oz+OJZn/rjfRCWv59ipRwOf4maf/MmQjJy1Yg+nepAUd+t44a
/OPvpqmMtt1iO5F2c8ptDuwh11YIsm0I6dRtEB5dklhbRLbgHzZWSrbGI6Lbz2K7QxP/441ZSb4x
sJc4rHVnNw2bSsktOVuGeK7zxXaVhijIF74fkFrevQbwS1Qr59XE2Ld7bPC+Ynpv3POZWHchGaY1
7yYFNbgmepuzyssq6d4ZadA0/8HjWJgnt/iqJs5Z8J1/dZo9V3OK/an+/jA9rpmpXDbhZtcDWiGk
AG3gYRZ2Pn6hFMxSRfPmVlRnO5uWDwlDxrjNAW1+N/NeH7PisbRHQzaR3DJIGPWTTfXnWUyl1TWa
SzcaCWYVhNhklh4wK/MVF0qf65FAALfmOG4l5uQ78WzkolhU5l9Mt7dgJqa3l0YoW78hYbR39qRK
4ujfINu3HKVsOlJL6nSQEf7SdxR4WgjVCsn0Pq2Ie0xT9Wex/fhWZ71i0nwz6B2zKLefJB+xvf5P
obOjdl5saHjuY0lPyveZtOdM/gP6mLMitqnAHNKSe+wj2q6tBIjU3w1Qg6dbTyaZxMSGFgQDofWS
y5cdT8GTy3LB9FiOQyUQiUCV1QzrK8KxzhsyG0+i0wfNB2Qb3BU6v0nS1me3b2nnthkVARKMqyA0
ifn1k7EJsRXEfj6rwJnkIVIyFX1K4LSh0wLmTXiCb1YWCMmTA7JnTb4xmpu8Y0HEG7b3taEj2vHm
Nw18FbP7JzDgexAGrgxUC/B2n39zM5fWYhuUIjExR9XJZIRsPEDlQbgDVYA4af9vGW32p2hdFX56
w8nKpifPRtau9hP2vUwohXsonTONCZM4DG1bfqegNB0sX8TVgOV0g4FFBxcqdhFVUAu4knbuLcyi
cBcEZ/Na3QmLAHd9RglFzSk+Zw2VRQVfBH3DL67KGdtl5XfuoDGuPpGieAj2r9YpiD7Apc4lAhSp
DgzXk7A3vPtVP9thCirzj2dxjOtD0hRF7f5VVSOCI3gxj1i8bzRtRTPP4f7JFtiykFWM6qT/61JX
tj2BE+JIQm/F7I89ysp3DZlFjQN+lRVF8hXu0XceSt/aEz9NxzpEWLdNF/Jem9c5+bboAY0iGupv
vuDAyt17Ix9/C8FExsRD3BhA3vigSttNQQXl1Dmqz9xEuGhg44MukRnYtG6d5WIgQDMIxNp/EDvX
egRvbq+cRDsU2hkze+oG0dWKMB1YrvL2Whw5825Oyp8ZXO0GNFHUHD3Nk4mCHRbLa5uXDOhjqhxF
5LdT5z6AR0D0aeAp3WQ9Ca2x8KwY5EBB6zaylmxSuIbJEmELEcsE5/xgxRU6a/D76gRLtMgzxn9p
27IoQkG3ENUBwLJXERcGRF4KF6HJ5wx7e7drJPUaLBI/iY6n7NxhWOxZ031o2TL04aOmdZOrElgK
T1OCETF1PjovU3IAddiU2JTGtM7lfZxYUhxgCmK/9tCKZHIRXCZQQPPxi4zFgWrSDJ542t6vQwZn
FhcD7dIoVUkVYIfdZknMw9pExU8OMJlq1ugERkMiceokXCOeSiWub3LwIGc5I+2f6gUfSi6fahVu
9vNUNdMdYRceM1vY1BZqJrqaZqQFN9/V+Jz04NgdoyRQ0wZJerQcjFZZ0eaX2g41KJ8TauduX0Cy
mtokW+dPydmzOLwMAnYxndcd/5MuWloN/M3UIM6hGAwpkQQlm8Qj/O/zFZ1zrb2XaKL0rrvgqXwP
BIAv/RZzaA4yYEFR9ydBcYCrEL2A8Z4s6ydpDrnz/E/VWeP8WDOSpreEtu/wAnpxN9pVVE0izok3
cE3gtyCH2LSufd/lqIbpBZlQgae5iRi0yH2I5eXW6HXXHrPnY0iS5mnLzj1gNIeqq+J6ywEunMt1
k4vIVgiSwP5YSbn6197EgFGkWpjvTch27WrrjXMO75i4vFuZ7K/4VSVPbrkNx7be3ipHTQzfl36t
l04xDi5jzmg3kx7qffo1YZ/0QjQMOqjobUFNC/8OhNMBPQLL3zfNXWjbkMp8LN5664aHUCDY/v4J
OoA4bjUigBT+xyShPWCbBLBgs4InZWmdIwstdgwPT3eFkBTan8fgR74ajmTTdKhhyNYS1bzM3y17
94xr1A2E+kK/oQOrrbYxFvZR6+dzZXFDHKCINPe4WDyYe/pR6znpgyTmbecm99ONrj8OomCfU25S
e+U/rc0x9IH+HdA8XiSZ0ENBzMKFZCkQtxejxPD8axeZyvmmhzfKQTlYCqZ9W8f+eqXu0RugnXsg
InmXgXTolhvyPq4+C4YPzJyCkrBRpaE4w9JbEQbI9EAXFNY4w4tZfNvGmSo8KQc9l3KNyxNxRuL3
Ov+Mdn0JDfVkcGimf70t35CMXFJVTu5Aaaj6VVoMhBTRTFGUIjpbplyR8rBaEJbadA0jF+cOJqEq
EYyvMz/5pu6MqQvo218tobQfV23msumoy4aNG2T+qjdL7iGCJHDLqx/et8xpSA1X1zj6z9wrZyHQ
jOEZpHfegtGQX0D9YAkTgAAA9YfLtVmh0HNKzS+xJ1f3saYecLPD8R5O1xdcal6c0G1Inuqx7IVs
nx2ttcxE3mCdM0aafqAj4C/TFBreBGWokfsEr1+WCD5CpA8ue3hvXuG1eq7tbY+EXr6RwWlKa8zF
o/w0j/XTNhMAH9LglvKIiWu9p3TdFaG6DOIa0sGXk6f1jY2b5AkjlUu7nGTJ0ejVjNp9LQA8QM78
dH+dZW8RJtJFUMNGfrGT+uK/pklKji6gjMcF791HQ10GJyB8aOPrzVlDKzDMsp76n+ejXeD2etfz
BBfcBH6GcOYtj9urWxyQI+GJHGn2Jwb7Qtezi1EoEe6X4ZJedHPOEaxVztVuEui8mh5pDcK+mGly
r7xXvqJEEF3asOEH3pvLJG/MSKMK/LsP7nSzOkw2qNANmvZ+udmOdzFyeMIS6V4YPjXnPWtXcKPC
wuUUI+gFJIcUmv1brvcjFW3B7/hKCMPOuNTXkd2Epdg+7GracjebPFxCYg8yTf6n6+w8GFL0uYal
9w+arM5iVz35iP5C2zYeRD+WDt0H2esgvgD87m0Hjbepj2HZKhJyf1HU0BQSsvAUbtnlphcPxNfn
c/bzJEPq7CQMWk/tX9RZ2/EiMS6UI2mwgS0FeQib6ENweg0iYvM7VEVhE9LIZMcQ4PXLwoL/pQGD
H/dU7DAC7RxyralkaxjFz0yEkTggts4xgiIZE3C0jvvf2FlJxI47e0f3DKlTH4lzRQGhwrFpRJg+
nc/1v4dU2N6ks1yOLGdqFHJEQEmvmP8dwZ4ZjXEY5qedA/dok/+JlwdEvjzF2DSkX3irjw5jqHLc
JwEUvSklcRbk3BX54nWXsxHDV6cQxm99824k6b4iOz75Q9a6Ndyah5G6wOSvDas2Bj+cK2vxht0Q
QgRbvixkBGH21jPGnSCafabyIr66DiMA5EvJbMTOWRzAqbsAPm4j3yTjCkaOFSi0nhZxNku14YKK
IvgJAxD05NIVdPTd6yTFexrqGkH92AXV+IbvqUL2JN7GTZ9vmqaYamNlTEEOnTqC3qjTXvBMDf7A
YjM+dnr8VfXQ5w5TOm39jZSx9Mh06rRJ3yBemUb1cpEbH9tsSrUPjd/1Sh/TVulD2vewNV9318E5
vtVKHWhRrJMbU5EedpoUypiMRnBQ6DOlPwSIRZ0XDLPBtMIMdonYI9bwf/KjI9zkZohA5q9SvlfV
4VQTn7BG6p6zfJzUCuk3LDBA8q0obs3sxN7vF9r5HTyd65Ei+Z+hPxuc9s2yio35Z3FfMlX8p/Oy
pH0ilPOiDDOaWlKC5YHq+z6QoDdFU9i7nif9bS3/5Q3g2qD106WcSLuF8eMl8PohSyj5svfUMx8f
bE5JHXCsQvLo+athXDJYSz7VX5RCU+yRu2zLZwPcOBTAKAa0x0T/3qTTEAKOqOvNJFSLemV3BPr+
MP7tKjZvx0Dt5kdAve3nYQnPIj+GKZ7PQh7a3pGs11aZTHAoPFhrIjh2ViceAv9Kaa3zZB9uBJfD
ox6PxhHkSD/tXMmzwXEc1TMwcFh3MHZvy8ExWHEV0++DstfsB+CXxlA0EM5mcQSgSd1hNSwJG2W/
1mEcUwJCdo0AuBZi/5do1KASnn9/szLCY+rBoc7cFUoscEH08s542hJCj+pUmZMI7m4aWPS11+vh
+F0EV95gQyvvtSMCDgM7Nzs9V3Dht0wUf3vmZnAV5ovHiDdoCtpPC9ljZ8Vslxz2nfW1fB0TJ8KN
piQa7L9hy9cNIr9HtPxUDZwqUJaD8c7W6bKI0u1As3LQ/JnNJS0CZN2Q7VAlBctPXO3jYd33y4bl
wO4xPX5tdCwrM2uJGIzFWf4vv/DW9pzb5pCMfPR+dEV74nCw2G2OPQSKXyG2owzGYEM2+up6JZAt
taezvGBhn65YBu72mgDy/0D83GtWmHKRzlmRq2tLYg2lU0YN05gHyDm2IMsA4G1oHov0puMFvo6H
KODzwTCSGqg8KeeYPIL0wIWaSDB6MO7adiDTQo3zALRwuhn66haB2LP0ttWj3joUDv4af7SggPcC
6zx0zpNv8at7Ge/a0XodI+8G73zK1GuHdnmqYFQe+qsvfxXJRUANzfunFTuYTYTDsXqTvD5CGYC2
DGDRtvy+oynxwjV6znziCEGhNjWt2vmxNS6LW8PRavxNAmZ+sI1w6DEX+S3ms0uMKQ8FRojUJrZT
h9A4DMDHmeniD4jbjV2rSMROVwdQWWXHRGbzk5EXJ83JfiHTpQPsgyPxn/sOw2XIGzG5HojAoLYv
K5+oy9khgBkGNZvPuK/1JJRvHRTFMjIgDqskvlMHi38Q2eFCl+3Wz6jZQpBhDuQih/0dQCikWWMf
ohOG0iC0hU8c/5sReO1uMFTS7xYrj6E1vOCPK1zmjzDHj9x83dH4CmuIm4HYwI3rLVG/EQRybwBT
IflF6oYU3XIizPKQM0m9JTAjqGOd8KU2Um0uK1o4yKCSejFmQVu4n364KFyM3ahjdvQRRKj6tWmS
Q7rulbV93+hBti2gsYs7RllG9LXcn1aNmBL5RdGKyLAABCK1pTKbUfxXUyNscpUdPtxZZAjzI/K8
fRvgd65UsVY4BaaUDl6xE6tUPt8i7OLDPHFlUo868cFILXZkEjwzIaf+9eAG29crvA/9kOkQKgY3
BmLkN0ejzjYbvleVfjQNryECLy+cLaKENXEsuMSyPHInhb/UPUQP/rRjF1osYs09rzL6b7YZ2E6P
Nf9LoPjlvJ1uh7OKNNauE/eWUgvJ+5QnERIZqfa6SGvcn834mqROItnDi6Vk0IwI/b+74+xCH2fI
BwQZcb/vzLHS7XalWa4iHQ+oK4dxWkP2SAWbm+8mp8uPUj2rUSh6UdT63j/3MnUtPsmej3tBhzBH
bekYyU0LAhnCpLL29ZOAj1D8NW39k54TGgN8Vor0ekQyYUQZEIQ4VzUOfGw839KO0MqftX88e45P
8RtIa4sgAKuAYZQcPVLhx4iF/nHCg49rDOC9O15cvk15sDWvRITDUgfYcoLSM5P1WvAO5WHFhjTY
x7TnIgAqH1GyI2L9e7nyj5FNrsy5Ux11yvAo/P1/v9x7e7bY5u1qlRk6I+s1hp858Urqg5dN+izn
0mHzDhFF1oa2d4lsJed/kl3Sw6euPKKN8ARcQSZkyn/wEKukLDppKFdIAO/ggg1E7VxmZmnaY5vV
3y1d8nGG4ENYwucGHciyM4OlP9JTC330b1nwefF4U8ArKCxTEDWa4twzqO5Wx5TXoWlXKu5YkOPD
SkN0IRxDWE/M1fFDGTY8Kps0jaZ8QJExy1UTSYM+0pETxEIIWq449O4jaR9J3fIl/qm6fPwtHPDm
DFhpkjpTLYF2PzywjdNMR71J5kXlWEUNvH31Z47rSZinHDY0puR6ig6cIQK2l/la46AgrsC27AxR
oZ3KwnR8M4GkCBSvCXbcAEvKm6A1WQNKL/d5s2VR9YzhOpwlnyHcBYy2Va4+1gSedzawB2LCYH3D
FjhOv1Ni7U1t64oxbDTFBxp8muYIA/RdAgQhmIvB83JZag+zzVaFgz5RNjgQSdXG4glyC6zs5h+C
MCqXupP8SngMeF01Te//jOeDf4Z6l05qXg0+D4wvev3e6tAsTFfEUf2z3AMPZir3Ox2XhPvSWeyz
EXWsn4QFcSiFrP+OtX+InvS0Z4hFhGv1j+yRVLY9d96pBEYrkbGcjtgXJV6hghEmw5/CHkJ/wGcE
ovp1QkMeB3n24ivmPkeRvvoeAukWlNOypIDL51zIEoH4uUJGmIC95yi00dUkTdLgQKRey5cmd9ph
3g3T0hGtPHlENXfGP26zuHuEiOyBEi9lB4JPtROnpgPWNs0elTXkN5PQFjJJS/2O2v1nB4oclT/y
lf2HRXGzgNOBkJccrdF2ny7se8o3/CAxCtd2d8yGOz6f1ymYcdhY3suwg2HuDB46sPZX7I0RHQDI
sblpEiPbTp3re2+vd1Hhh1IO37AkwVkL2SzgjzCRP2oE96d2dKsVfZcSHeHFZl9JA/jys3K1EdHT
n4TzMeMJjzeQkvIEs70cpl47YX+xNajJuzDH5ha/Hf15FCxAo0Ys1fZq/tcsbQJ8yTh+G+TgMn7k
bDukWfllDqLXXMWqHgKdqNTqJ1HTGFxnpcMPvsaUvAQ0fcVBuJYOIBSomvit4Y7JRfeelvfIFzAP
TD5z1VcF//KLqs1xNthbT4oyqmMGlBCZ828MfG/ExSZ1xO6diXEnsS2J9Im1+mo+PkTh3EUwKYSW
MN3Iqr/TViMwRgurKuLJtIbPtdhCllTffiYxWQ0s65e+mtl3UEEfm1fBj/yh8cOo/Zlz5lLCkqKv
AK5lFvZmqgwokG+ij7LKoxWcMuFJt0mfX9BCYv2cZW0FnFICF6HPANV32lYozBnJtN8XSYGwJiGw
OoNzdwL4CGwCxWJlvuoiZdQZN3iMnwNJIjY4jhJdVsK0BdsIRpQ7StC/+JkOPLgcMw0eVF4nmDTz
b4yxTL+Q/L/0Gdv+xzr4O0uDR7z4p3RBNJjstfwVwNBGy+09kffQO+lhSx+OJ2CzbkYwlazGK2ag
7vuuO7fGbHMxAr1fXujhCWmTf2z10GEeqUfBmFdGvNSbmuPLCGPXfv2HPcUw5H/nRnG0E/82qdyu
dgeskifWaPbxxQVLiGIa6iamHlBLKUqtlkiWWyAXjsvFMYCpo1PvxUWIiUQkaWkF1mzhwDhZwXmg
mN6wZnkSzW1kIiV62gSE11DFhhbg5+RxHenIej/XAsedXm3HKsjMu3Vgd6a6j5Aw0fDMD5PhhThG
AwQ5Vs67yh1aWOyD8Hzz+S50enTTjO60WKtBFGpG0wKJkTTg9czQNVca8fmGbCXo7BV27I8LlhNe
nGfA2/SjcnMY9r+ETYRQwd6x14Jwf0+KxKpHTYmOtlxE49khONd2hV52VwXcJ0laD63TFpbtoUHN
gLvZMFJFX4VvazgkC1y7LljDER7qsPJ7n8vRRbAR7990qDPL8DyQKkp6ibyrn1Vm4ltQcbtzgwaD
3o08sbnFlItChMb7AwolLDaBa8G1FtTrWGfrt/HXS7/32NPt20+MyILKljp9wObRsrvO5/WzPpqQ
DWN3cB8BdLXLLpdBXGWqikgNrshptJNGY5H3zAkIjYu8SskIHSJDy3XPxL+2dcEwUpkO/NblE4hO
FqM8P9J4Fqyf/J1tpEotYUpA2uxxoFDp5qhS+1WB8eKI3D5/qWs+sLO6k7ul9PmiVmd4sDm5HqAz
KvDsl9tWgJx+hzA8HjL7FL1iCh7iKtL0OgzsRiYGrtUHYtnHpZ1R5Jh5E97Jx9rbG3ehaCDkHSJd
IJlnD00FiM0jJldfow39MYl2/mPROH46d4D81vWySqGlNkNvZh8oHt08rrOueu2Ych1T1/TCCJI6
x9YMXJi31xbIq9rE4SSYerWlGUDoJ7H2Nl9Rms5rywG0/TZvCyP0i1GwH2NFe2qrFUYyPA5KQIlP
f2/0/N4uUHs2ID0XcMiWZI7LhVXHNJJ28EpG0FchFAJMMg5TZdQHK5sBMVyIrg+SX43cgjBUso/b
FRi2+Y06rSy3to0DVDnZr7RTB2tnLUxSHeZHvKR3aoGdZH0gMDYgfM+E//PS4Rm+947Ura1N6jvd
7jJK3R5kf5ozkrV+qNsL1m/un6gygDf7Z89BV9fLtdD8U6w6LHkJbPttClhNPeOJqSuAKwStmW0U
ZC8m6lULfU9Xhjk0yPe2yNMhGuvK+fKa9OLcJnFHUnwJEyom/grkBy66xj8ORoWhEk2LhnHX1v8L
CVUZFkCMXn948m7xSASEh/xufnormQwsNgEqRIMYPSBg6wROeqPtLU9/cp3OwJvwF8+YkdHZ3rAF
pKGphlkEFaQr89dtPRBaAHOl+4ADxUKwZMIu+STVS38dONzBN2hqx64TWLOS0LB240yfyzKdv1+I
nMvenWuPvaqD+PzPp/l9XlCbwqIfpWXwhKD9BG4u5Fy6TpC4B8TMWdi8p7i9icdi38WxVwGDwQQD
9zg7/U6bpRndIUYwGSCir5kN6alopICJtZA8eXocfpx26y8VqZ7zkU4JciUniu7wEpdKYxN3wKUi
cbGEwmq2TQgz/9WYBhVeMIGR4S7hJ/mO7GUCS1kGkKb9TUxh5auKbOpO1kQyXuDvNJ+Oc6tcb/lR
Xle7lzOzl0Pcf8S/91DJj4V0c/DMmbyVDID2KT0xTXvvhH/43qM70SN45lqvmnR4DYf9TCnkJnNi
jZBZsSURAmfOs9o77Nk/+lUUYdTi94OKJd9WDrk8INUJrDiu39QtRVPFpKZM4/r5Hdf81rBmlvCL
6rWS2av27jTXBwuJ9SUDa6uVFpt8G17Tb1Ugx12g/FkiXY+G/fqKNJrvtP5gLE5L2O3sD9R0mHv1
raTi3AICHkux7xqxyXKJ3rxgevVvFNFEEsgkyp1La3iBDlSfVg8Hu6I2p8SWgSLzXFy5ziNdaY25
H0rKgDWbrRzzd9yQ3dxpVdbG0NRZjhVTkzV4L+uAOPWBDmOA4rYNRwpfrsTefhnpVaZ0Ll/vZQ/6
qrfxwLAAVwwa/b8422jhqknGJoO9SXW4nLR/TWMvhCmpN0UZGTH6DEBn6+vwgYDQnNgRFv8KsgWi
v0nuDP6+o3sGqFSyqZ6y2CwRzcXZm+IAsYA9e/396OXwXtYl9dRQz9Vmd0mqNVKJUdeiNRnzYeDN
tAmbC/s/j8rD8sc6fnj4mGb9OJTYoXezOvTaTrfxCdwARpnXko6cZ5VWwST1+EShfDH7igfpdmOq
ae2kCJmOE5uVzNwcZVbXkUS/5nPWigzB/t2xuHeRr2stlw7ihNroiMFy6m2mkIwJJDODK+6oy1mF
W9k/y07NJIpJcgbEmt7MJUg9AILNoo1CDEJAu8xAc10ywn67pV3Rv2cdgDeAn3BecHp6DTAi1198
q2RtA7dZJRI15hf8u6AZAnN2DZxPsJ3tNbypGNHqhs/PvKdkZPGHFsVwrGSJV7xd+4+DijmgEZHz
S96rpaDyFRqEMuChVuVq/1qjeV3uUVAr4/K9dQ5m7Y+MUAO2u2/YdI/MwRNKumYdqIedApJ+F/j2
KmdbLXR//hJd+3uL7xDSQMeXBs9DIw8QOtM3m+MnmTeTfqTX/jWT77/GAACwyCZPdEE8zrXj3Pk1
+L0zEEqnjpffAEddO1eTi6QxqVPXVXofOFgn5k3zv7NwkKlN2UlDUz4J2jgkYVMuNAqx9dBH6NkP
cc549x0w5xmbR788njGdQD5WOwBB9wF6mfRrCFndvOgkpUR1+EYdTtTeCKdb6P6JH1uCFlouXDj5
yO1i99E1CN0FJPcvzOUY47g2eTZGXLCOQRuRbe/ciJJHTx1/7xLCpQMUMxICFAFUetj2spahc43l
XAfKYye2NRYJfc4pmPzWkHoxYKSQqiL6JNddOtG3q17gQu2vNSuTqfWHsa5GeZggPwJszOIDjvlh
Q7q7He7csvMQpjIZ6dEsZltjv9vqU89kA27R416MbIDS2IKfDOC3JSmf6mR6wLr3ogBJ1Tq0PR/7
/y64xxQuYi6AeYJis3nO1YSNr3E4hB8plEZoBmz8hWCCc1BMc05lKU3E24nNDwqWYJ7RWkSjWyHh
qX2oxVL+QSJTMoZEeAlMKb9M+3e4/F9Nr1Gfv/qyLLA22Yucekp9OltbkUUPVPGue/DOTI5zQmoJ
IMINNOFJ4FRZ6oHtl79uNKNIZuz+1ctyVyCupCiNcJ9v2Lwof2BoEfVE/4yMVfTG/VSezVOxJg0u
iRFuGSQ/9C+waxMi/Py6u4Y29FvaOuL+3tTg1iLu1FQSHB2J3c7zVEPMpU7l3xvfjEHa9bCXy+bL
l+0jVKe6dI6If8kB7/omUkpI4gQHdfOibQ5wtuaQb7FnStPHS6A1tkZbpG+sF88+OUM9ZR4HkDX+
ZZZ7vFQXtISaZdbUjuo8XDQOtWTmL/bnnih4AKbpCpfcYg+sk4hXcOKquuReX5vV3U/09C0V7VRQ
oA0VyjF5yccCMnf59eJeNp0uV6elmcwvruPKUZpv9mqjbjj8v/tvRfeMtcZt4XU8L3l42tJ3yygH
GLgM4z19zKtKm5e2C8fDCxDFXoZAlxShXxqCP65yFqpaTbvXPZxxyo24UQMCgGLk4W2r8yGvPPjr
OhtZdyuJR13RH1O5uIGdZnAZ0U/b13Mj6Kuw/ULvP8aHTe7NaWW/sfbqqfA9a1f0j7SdANeU8MCH
PXszeAElO9DL/G41LjQ943BzgwxVgIf3U0Ngewpr4Z/znc3VS+FUHspjTXjg2GwZOTyX4szdkrGK
uFDm2TC1zk9+qdywypjF29A27w1ZfZY816TnjWGl1cKaSDSIaJISl3j0ehDeRSuFUBCizt0AdGdf
dvHmg3+zhyK8TfPWvW4/2FTQxGeKZTYsB0PMnlOG2+hTp5haMgBdhYoiTAM7qHTOxZv7ZngIXQ8J
xrvQIMfPFOAjY4a9zWHquAN0vU9z1rZa3t8kncXRTX1Uxb2P+2jtK2B0PU5DTQv0hgPnOT1BENym
9HeQB9CeX0euTLilAxEbLDtRr/aLGKa7QGD2Nyic+g5jczFkftVthJVTiagTRlexjMqFMTv6+kcq
O1tifGyslGfJy1Pmgw2LpRKjvr2oBiJLrQbNLcUxe25sO2mFsZRKrMklM/35XYpyUbAi0Oy5Vgiu
PzqdM9xDdIxotPby3a/fMbmrI8uhkM9SH9p8gzdG/hwJvJW3FXht0u1AF9PVZmswruanONlFaegm
ZuRmUkW1ELAwFhAPWdj56/oYQytr38JGEZOEhmRV3hPMq/Uw/qN8OYQYfJI9vPXAf5S3hI58IseQ
1cQ+Bc8OIsEbC8xbecLpjpWw4kMIoaBBDOGHyW7ZnX8cSWdWMcNfmrtCi5Eq2LVyAE5aia0UQfkR
6ECGzQpiwX/8ClGqbssGqZ0u4+itdZXfVKJVWNjER2Bow9rr/hsbfSDx2QOj5oKSu8G/z2IysjaS
evrPhQ3ekoyuWRrrgphxRQFFGMXyT4lp3bSizUrpFNTybrqr6OKwOTR1bT4/WemnwH8pyDsBIYUP
XOn2+UYTIxH7BOInd8LaTtkB2K5Um/I3IQCTwBhWB5f5lOh62T2US/T1z4CibxTgFjJt3NxVhplc
Mtnx4BDZrWypk2qkE4ENLEt48sXRrQV1w7986nFg2XyKxwN4RnobhrXO6uHtMaLZwp1HMoX7RleX
B1G33EdcM2lnRO9AaHhL6HquTuQT1LAhldPVnOZgTqDIpBZHlVutZ5Dl4bvDArGnDOCGpdmqhJiU
QmCIFyzNRzIv55uFNBx4sHtIAdlCXdvRHRfGIDYN+bwOr6adeDISDn2lRwDGXGpRfM0PMci6VCTI
TTgox1lPo+WdQgJoUcL2A8IjDCc4Nnc+zg3SS67fQWU749MUo8M7L9eHd5BvcblhZzbMEQOTFItR
lLAw0oKPbSk4n+VYASpOLCfxjI35aumN+rc3JGzMZSihSMoDbl45VwD/xUwAqelZyc9jPAZkQZKi
SIe4AXeQ6RziO0AEO0PNW6OVo1Ro5pB8MUoSGe1UhK7UlW65rxSeP684d496TeoInFEHMYzdv8xs
ReopeqC/i5EgggdeDkmyhCVdXaW15tj+o4jMtRVVCSQrzxbCVrEYiY+n6TnWMAl1bjyGpWi2ZKQp
C7BUkVsnB64nUXPzqyGTBeu1PQ/hbllnh4gr5/fnTTSh+YDY1IqoQqGwy9RlVuQ23HNHeCw8Ffer
MN7X+kxRRJNC4U2W0AjEpy3u6ANuBUkMn/UVUUdKfFeZCVa4xqrzgEcCZyxlEG2IKQVuZVaESwTg
CeZChJG0s8RakXJxJSduwT89KTcqYUxQ9Kmn0oJwc3xIcdGISCs4NPTbT8/zWQvHNn9rzPknfldq
mGtZlDg1UgruvFkW2VOjJWqMCxTUtZegerjXyrBKXqtXHYeA2lHwHdrnIJ4GBieYeBMq1m8c5GMV
5zFQIMWPTJURxbRDDb+b1NRbRirzrbT5M3PNhv8c3EEzYGq4ekzT+Ydk5m3vjgl3TOzRZDHYeLeq
53jJhiSoCTEpI/qlo2G8SkfsNCcXr+oWYuAOSNuyawTtqIAoY9o3yR050eiRfrbj85vbrGyoFWG0
ETdyEiNe/Bdb700C9Gf1+aEUrfhC2/IRjsrRce2FwCDcobcCg7VTHn0fWdEWW9YUgPWLVVCU+Gow
dtotOqWOpr0tNMxvCJtrCwxf97Us6YdmrhBiX4dscn5QDHhTpGpMErOEH2HSzGG+zROLhBWCUe2A
66kFEO7+17oh3VBwhpzkGLSN4foy2DxEbGPsujpN7jI5qeGXKeOypGGhjoPhW146IdhUK6oJVzl9
bgyAmR9gdqKKD44nykCqHCW4OoSc7P61haSdD2xDkDpA1PSRZqapW62yz66D/OtK9q1+oxpdZ1cV
EVxBSPg5G0O5rcfI7AMna1dQELDiMKuxaRp4+b0ii7cZcyHHZt1B8M6hFAVRogQmbFIIj2qCnbcK
jpWv4P+WMtCrPu5HHdizussud22FdEPCps1dSEzHs/czxl1dmtY/T5k7KSiS+azZ3c0fCO/qb+UP
N5fhNI0qDTUTppXWSk6riFreGeA4WGYUdQaIOQlhze9TLCiOu8guRSGfW8CzZmZQe+QEcNt/q+z3
R+Ic81vJAB+gWdua1+YzehNblBHmNmrWadHbgB/J9tl+WK00cleeXMhZtzDR3eaQbGNjW1jAlnmZ
kLeSOCtUtJUUrJV8AOmemG24sWe5kzZncqvY5+92gL7tQe5P0O6pbwqEayAUxELDi0dot/56g/i8
E8grMdnAJ4/C0caBjtGjklPelgS2GEU6o7F+vmWYd4omvAg8QHnkqO6iDWp5IGpJil9oxRp7vD58
k5QPwQuz4QR8qjWpqkjIrgr6dqaz5hrGSA/OZwjaO2R6VMnB3cYTEToZ8ylBjaCH9WviDdRMhuRq
vixD1dIpHN7yQlduNDwNUdaAYRJmo6aAl8YH+pDafmm5zw4lV8ND/T/F5+RyUVIjTfljiLIS4LmD
gWlppHmIfRTXm1xNMxzcu6lRjPb8FLrUQEYAhyMuBefKr8qYrffSlLrgPQ3WeHiWOl9gi7xEy+8w
nX0T2GmLNN9RiUk6i0vVgNKP9LnZtcrtg570Uk4pZ+ozF62nMOLczCwpU6uM+vo4OvhMXDGiDBqf
4APax+AC9TKALw29zodAIp+Yi8x7BByp61+2kzEXw3SMGI53hE2DwGyGfiwFNH8rfn/j6PPAluRF
6r77p3RD0gKNPtSCOnEHp657RXPmRRQOdPevGwyY8kVEg1tdgxrOk7YNJP4HbMreApgrMr2AJ9og
B2h3CL8k+4Fq1Clr/IyMI2Kq9xZ5rWCqO0fGRgpixxlyccluHW9/Nqi5rhMwjFH4XkYuLIBw9kjE
K2NE05MJOGY/PUD26QkDZqqsRU2gwW9aLW+1nOjLBJusWVs6isUYs+Qvm1nw79+aTtC19tK+T7Eq
mciNe83cL63ELyVJR2JcrdMwOqB22hEy8VDjvVJpRZdcdBIg9Zs+WrefacX5tsBS9zo9JdXR2rB3
gM8qMTdiXk4qWj9/ru1vAsHr6PG0kKpuCFr+AbQXl/d3saUEet/FaI2gw8KS7Lm6CAOxvann+Ifv
OJDwdJXWjR3h3R7eQ9M7oGkzGA7UcdK3Lsw8qygwCwLSLZRvoHs7OEX+gSNMYq0uAN1kMrx9wPQy
eJKI278AtXf9CEbSzVYDXITJyWjFmAn0WPHDG811JSk0fW8syZmzqNirTdrbw2t+J3lxxT6gclAl
3dEDuguUpF1HcQ1uehW4H7WMk0U+8Yk9uBovvELUewFtL++k0EBqpVXsbg87R/AMyrcH1AoIKnQU
e1TiVrB9gmoj8o8uTXyP0sY4wauc3PsRv/Ri5rXAL5tKFc6+tfhhBk3eCjOuSBSWWjJS65vRY5/h
UYU6rqe09VuRH5Yxg1cCxpCHNJlo1/GmCVoyKvzDc/uoEDdqLF1rP9aprPB3/3fZCIPXZMcN5DZ6
A+82ufI86fuC/NPVOOx2l7IDroA78VXi6ut2zDO1Sky53PVeOo/EJywHLf0E6aAMQszee6s2Q6qc
4vf0gpQqP2qWVBiLlhbN/PMhlJIc1A+f6qDqD/JmYlT7PtIkb54cbkGjyOt9tD9hWe2PYurb90qW
ta+M6iKC9pgzIEeUfRgqo3l0ns8RkeMrjrhrB2OOo1+3jRTzGFsER2xh108jUcH7TbG4v8hBhzEQ
yhBHObMdvxoaBy5CjAL3S9WfGqHOAxYh2gDujy5O/P3cL0mWIlhd2fq/FQW8KwOayK7l6yoWeFqq
1YPpERTDIdiPl/IDABAiq5gy6DxZ0kz2ms4rg1rgoTv1sUBGpGncQFRDBLHp1ACxG9z8vi4G/Ovc
tIkKvCidViIPi9rU2G9bb9QMrjps9zxIZTDeiLQREq/txu7b0bsEW+8gK20pkMzaCwiVfGwY5oiY
BzQsZj3ouquBQnYBB709XJYqjeBxdPh5Fhl72yR2RC/WTdm95AuCVr+MYh4X53SETta7LJpCdVUJ
EYmhnln/CJ8AzHQyVxdcECJ67QLNhIvKzDliT/BuJ0IfIliCp6++XqXmsK5IufbWWZkHCew1azVY
ZCzcotcZ1WBEzefR3HZDll+edXkQhAmMx72X7567DlbPUNwIvu0a6ePTl9NtGKWNDRbjn6S5X544
H9T0XPfNMYrVJW5St/FgHFhG2xGknB0iH8q5QAursrE6Y5bS3k+5/3OktLbn9btjhyHp+MAt0lJn
rXlPoTRFaUu8CX7oA5O2Yubf9rcs+6k/xF0HkDJcrJIJlX42sjlV4Xbi8Ige3TSDMUyw9w2CND1h
3ghYZsTEBkWS/zRauihp5/Pp0rvaUr981DQJmSA953mxblaPSd1UpmRUM/bqXi+eyrgHrRvVVLhE
lwoG1kzvJ8bdJ8hZE6QJAHztlFZ2V3s9f5PtsWEVIpIUP8x6xnDajhKshQlVSTvaPeIBORSn4/Yr
BJDwgNDFucLXQUCDZOkpIfgNjHg1oc8am9caL4nlmKObDPvkxfszAIyDGSgxx4i0Afia6/sfEWHH
axB5d0Ewx/Y13tBAp161m1wjtZs15dro9jn1jUV5PHCW3CUJV+QnQydmcQkleX/wM1MSCoZh+uJy
e0kcXcCer3eRfF+Shheun5yiRk62viJuWtXigArD9Eh3EPy7rKN9UtR5CvInrDtQBF4sInQM9u57
nAOG7yc2iDEeebE8nI64N6bRMzv1wnc7W6RgUQRz4Wqiddkgo0kDWRfqSUPUdh7AT785GfG9ZQob
P8oDOsFPYT8964CBhdg5M/O8ZCSh6YPG6DcoipZ3xgaVMz2nWM6hLmD1butntyUVWuNq5QdDqzfz
Ju/WIEEFOy3/eJLYk3tkt9JuqNUmCKp1Y4GVDmNVk1Hj9oURln4lvKd4VsJww1eEkZw8ns6TeaWW
dFIfsT8fxgBxCpnYH+SaTQTaJfT5wHERI7SEMUTw4EiTofwh80ixHSI5JDs/fADchMu5GjVLjjl5
GsYAE3cMWsEKlC5RgN+8BIMyJlDQ4DPK4duvYdvOR2SNuDaaM/Cbnk6s/tJljDurj4sof0EsGIGd
qxFFOCvhgIcvTU0Yg6Pfen2UwqC1m3iBaz0mjbrKuAO90H4qzXMqmOPzSsAojam8lGn+HVKyygAh
4oZtnlSTF0jN+tgkc/UlxHbWYrKD/js8ezv793H6oYI+x96pKRH8I96xhajAN7gqgWA/jLCMVCgq
H0yPZzgebs5/PXKHzOXc9kYCnbItzyw8UoNxKSMGBoyBnyYPA2QPzDswy9JiXBsHGYLTYScfCCeZ
Ox1RwxkWzJdQo6xf6RPpoW0KGDrGk6IOyWlyXSpyjVTVKkgG3Bh9L+OMyg/M2dBegPYHcejb/UL9
E3WSOzIvx4xku5PjB9gvSN+LXkl3BojDuJbrYAzR9ikeffWbNlomrZcuzWFQNvuPdv2wRCrtDDRx
HD5+Szw9xJ91i+nwu43L864QMF/rhpw6c6VwRCXN2dg8SrXHpSdwgYLTvn/Z69w2Qe9LM/EZ/2Eq
7xmOrfUWYwjFo1jEQD3gndsThqKvFjm3al417PBtzlS5jtOjpWve74kkfQd3URLI0EE8FzKcFI6J
COwxzdEApHSVr9leRfgJBAdzGC8HisAi9xVc4NJfCxRpBWIrFY0sXf+xbE/xq74Ujb6lQcVSbuOW
NUlVM9MgvAxjRnN5b2hGh6ZYT6z0Ps6HFte7vJJey+5IKBDeYPI8cmhzQIKeRnuB4Whbw7eys2mK
a6WfOAgbzWpZgnIw3VRG1bfXUySywvF0yW6l7O7oSRFotg+xBiHt+vzqnCwNZR4pJznJKkEGrXfA
MVC7+4hvH2qlNtu/O9h/d0OpnNTP+5U9NX2dzXYxQjHbB9bjMuUwWX3frQlwJivRJwylzwhbR7RZ
/xy2IYzxLuqVhXFxNxr9WpCYm9rHM3ycavtoZTlJ6yaWcpysEwerFBdPZVzeTgR0RIyis+Hg1icv
sJj7XgXT8CGNNvTb0VCaX9vFHsG+1WnaTFlfyEPR7Yr0AQC4215uvM+TroVLNoWpLquMX0XCoy3e
tCxa/VCAJX+rjRzjqFZg8rVUhvpZ7fGqQEMTppf8CG6o0npv/6Nrm8wEmdpVCUAp7gj6WzjBCBw3
Dy6/1hCQIMuJVmff7M10T2lc/VAOwsO/nyN4DcBkQzlNciRAZsh6dEdR2qUxloC2531w6YY7spfC
ITEMKu3BLznoTIcpmvGM3AlELPMK10VI8haz7RIavMsoPEWuSOuvUlvTS3l3LKiRuGgJjozCCyhE
MoGLma9ilaLgjLxzO+nKuLrcrWmqn308Kmmpk96/A+WWlowLlrqcvpR1bFQk9msPAshO8jYtv9iU
pap04Y42JUFXzOSQ0NpgS6wKGdxVCLCJbOAdrmLyGx4NZ7E5ZnrR1CLWELEWsg8q3K6FTX4lBFLF
081dvWdFFS0i+TjKlGNr+lXlNOsbTRTFMz5XhgjChWPTMF1tFpI87Fw6n67dKx30B8U6FO1GtWm2
0dGVzXl8KIJsikHEGAcv+Oj/8WfWfpK9jzQ15gE2M+9Ig883+sT76MAfIAr4hoAC4DXkjqPZm9ae
s9xX0nLiLxpGIUEAt1Vj0IgGT9DjaCwrZ/Awi0nWcDjh7BcxFa/kV7IrTKdNvLVmusvP19HOqgK3
YxDLIEkuL74U3xQ5HVzlj5oydmj3zkWohC7jfSAJoZ1AX2UNYEMwWR8a2dXOOqFz06VzA+m+aKZy
3Io5C9mPYZvEeIyqkNyEu8AWSTYdArIDDvK4HFusvXAYd91T3oGv6X/23MR9adhCsm0uGIBKDqXb
zbj+tSqwjrPWH0PQPzx/rvGqPDAl2QJbUW8u8p7yF/Xd3b8o88/B84zP+aZyJJ6rj9raCgZnu8V3
Yzeplw63lczRULXjb1cuUXi18w8bIVqM65MteCLPjmcfinXOSXbK8Sv3mwUVOI4sNO4cf9WcXoyS
EqLZ3ZzdcF/iI+871swCUEpaAiBWcRS8sHZpDhhcliGHtuHrVSubhx84ubqV76p/ND4Xyy/lJ2oT
VE7FV9aAN1NkHAQ9AHCrXEFXIeBu1oMvHVOCwxz7bTSB1jT+BdVdNNogNnLvA/WPQpzx3cyJ4e5R
JK7ay3ZPKsDn+1zdxOWj9Vrpi60OfXj/H3/rE3SdJoNV/MojZMO3VXbCyNUKx8bLGg73+mGTQZEJ
CxyQL+ZCAil1d4K+dwtYNSIdgUGdNV8oXeB4LfI2oZsFeFUQuLVWHL/+sRDey9O9dw6O7SjaFqu3
PHZeYx1iCyXXzw3Pux1IBp/Yx441yYzfGMMBQGT0nUFoVzKf/bhDjMWUWoKu0NzVSZGoyN7stKWL
6rixkzoQFj3E/RTSQeur/P3XNG0KggWD5ouoHHDVyLwnqp6eoxvbyuoj+zhiNQ1Bxj9mLgvIggQs
ydA4muxRFymC/7HLhEyVBzM+6vMdM4Zp3GiNLILqWeKi2eLX+ekSDP8334pab51kZkv6ISlBOw34
95qPFKwVmgi4qXFkn5iB8NWgYMHiyVcgWD37QEuzqZJC1wmW5kcUh5egPG5ywd62bC6vyWqYqPx8
jFMnpbd4QjrRy6nuEQshxyt2bhX2htRzCNIcwZvvqIPmyRq5XPfWiueNOF/vd1ctey72h9sRk8Up
9gD5wp2dLJ9eLM9Q62Mm+9ylHbVUKcSnssIZxFIWldt26jGnfAq9EwYpor0n3bxCvGhfxn/KPgn2
v4gvBIMZQ+3mPbar2ZPvj1VYTYR5W24L10MeJKqxH5mLpZSR2V7JKG4IQsxp55k2u8nnW4u95VUi
14giTrRsXtR4ylMcpj/OwxjSvOfaj6TwLD86khtbpteqeZK7GqBLpXNxs7LYu3/DmCum/w3Eb72i
j3jws0wvLZTeYv2JdAWbDnSHXe22ksYig8g/aqOWFXISFY6BpWCDVfpTRcEuIhXYAWXDOm+rDTE2
aGrqfgW3mA3xMk54+FUGC2Co3/1SKuB+37FEXnmLgs3nNk27u8GvUHHZmeu4KiKeIya3fEcqkGIB
e5Kf6F6BOcKm63NqNGZTLDFXmcN0TuO2RZCQkAO++/gN13oveqbthTomYR+cxAxXI6/pmfS1S7FB
8zusAjwDDbipfes69x01UqDNwTQCUvSkMs0lske/3nGIBxCooS04dUexaMzSr7Kwi9rvRAQKEQdn
QHshxD3mqxlwgMEhpwRY69RvHa9Pig07VY3oVT8Ns/l+bBd2XKTqXef8+cR54ROmicN7yBlYSa2+
blQ+kDhT3HXu3czPwMj4HU/KjEugnzjGBeqm0MxnWQ4NfqCHBblXAdE2JvXWHruhg1Vxv3sTxhYJ
RB6ybJGudyGs9M7MjTGSPxfF+HA/Y2OteLJr0PqsPjCz13+XkwKPsK1M+Yj3DgbIokjibR0MZiwq
HVhfb/vguODi2X0DfyLgu31iittrArvoRITvcMPbT9UNq8ry+7Qg3CsnjWbJIk/E2BpVUvYHhSuU
D2SuPIaJ+F8xcyL9+jv5VeiukXyLe7FhGjmkcW7we5W4IaBemBbmNgcriXuUcKUIiMOgXDrixB3I
LDU0qwk3WZiree6AR5ddPCKV3zqe2ZX8k/9Za7IDdYugXskJoJw9jsEFUu44m7wA9GBdgR4hsF7d
lo6j6z3wbqsDLzCtYEkZY04eJ1V3Vr/SqVpImSdN/RS/sj3G15xEws/e0eoaFTc4aVZ3TSzO70Qu
4sWVFEzAp1L8637pL7Y1COx1zVmvI5Xg2KqV7RnSBg7pbyq6eJsj96nQ1iyOmqkXhLMnM748SGCW
W5qR3KElYKHOAb9tyjDdiwHvcw9S/7uStNEU8inD2FTPJ6ROTZz9z9CgQxdSTTpID2bkWFVNLdn7
8AH/C6suJu0wtITWR9/DMuftUK6W1fM94sPtIoqlmyLhYgL4WSEcPWdHno8MVlxuDoFPQnc060ch
aDNHRr2Lo9GUs0UaHyzdw27vP7DU2GabuReAJKqHSnsThBFVOHnCoDooBqSI48l3aVvKq7QdWo8R
51qawgRhNKp1rSNOZmyFLKl7HLzuGRdftrUKG/Quv3RyUtAnaM40T3hnLVhtJCXjsryRER4YcBZf
oBdZL3nyEUIYSvhJ9LrYz3UE7NBDdZOwaMyiwrPHJp/aBIfQqsHyEb78GPAm+JlF9wAQi1pUEv15
1lCSt54fl+CWq3824e9zOEl/rUX0J21ZqveA2Y0uPXSO+YUgZEpPC1fKBFHy0bsRM8Z4BMKCqsam
prA73EO6us4MXwtCOfs5HDl/Fddv6GE93ezW2O1PTARE7Ubf1BZbaYzTPQ3b5+yT4tzrv14PeCzM
ds0Qo717H9tamuv/GXNCBfO3lm/b0Svu3rBXEQUBoN9hw8sya0x1d7lnkSaTq1UHs9KiU38Ov7Yl
6rw2YuBYnBu37T+9hQSNFMaGOe4NazQ9fZ9GXQZv/01caMdG1FEcloJSg4N+m1d5wUgzZU4PpX+J
cb/jCWH8Cig3yfjvtpoUW21rsReEtYRjktmiqXmVrQInVCiESjRdEmUze0t2Pyh8XFQlxrrzOAjd
HHH214kfGFcb8DdjZzodDoVORYVQ+eMrTIHEUnhEGSCjjiFveBFLN4QFLP30WBDGHAdZGW3V60H+
D62OttjooRr7p5jNAXT9Qaztoe5GEHaBClPaWVcYmD9m8M9N5W7Tq0mY3a+eK1n8FWYip6SKHctQ
UUM9KU/KvLpozYMNEI5o8lN1UGsJU+thP2nUAlQ3Cy0RboHiQQx7DSx86IvjZtlgpKv0HM4Vf7Pm
7z4MZkWjaCl06A38xH/Hy4AInN+U1zMq4qseB9gA88JfXimiAgSN0hQ4+0qTKcxDQRgP6AdQOqh8
JaHVF8paYKTG2zbw08LcTvMK/FpemCqdWXKcK/PyF0HCzQqrBiKn3JB5j11s+lymYcHz38mI7sPH
MQ4PHjVqsFbXWcN8vmQdWMxoonKrAqkxVWWnwPcFfRsAIli4wc2tW7pxbFfcnr7vtHPfzb6RxbI0
o5YKD0luM3dzc/H5JjEOizDvCezBRGwwH+DSiMIAkO5OFlzKC259OuRpf61TjSAMlAxavuWOiTFz
0zEaBhQ1rod/pxecA0WNywzmBTLzP1r1MC3rOPHIodJLCF6zcVSE+Z+oNK0531QGgZwhXP2lTyno
R+hSK36qkPm7pCFB85KhhAruB57RTA7s7Hcmt/0i2IfYAWT9+ZUTqWf0wvLxBRMOEw0aqqk9LES+
C4OkOnEMlK6Vq/dh22tlepo8dlr4E5W3fo0LhoNy/bGTvXajXq6Blg906mcTjHlzV1QfzpdripXg
tXHvNivXXyfqRs3ZsGybX2eu++oR0+TnkD2dzpp27eWV2Sqc7H8V0WrQVW3nbrXg/TjjUcBYDCoq
lilV/QbQazX9kuZcwN3IgIgtDQH+QdPsruMl/FuxgIsl3BrBjuWXosquTz8FhVeqsbZs/K4a5ujz
+e6lnFfm1Nk2CNowV/HNzo2G5Boq0PjD7ktiWPCWTaV14hpiy6BKjAfAku7VTXpU6IrbcuX0Pw5Y
K9SOYXrRyQaNQXyaqvVDXI7mO6QL6+hZ27hfV/mQ2SJrr7KOyUC1GPNvJEUlgbDno9dfQqYk9BoO
DxEIxNY9cluSYmjaRrLwFh9H3jOdsZ78F+9yW8/ZxUCa6KTBCwoWRUKVN9f4w+d+T9jCZMxThHrp
on4IjuyATQvFxkMINVC6HldaU/wD0vWuEjTZ3dkGpykMWZmUx0m7t6rUoiqCApuO5inCL5b9f+sn
aN7m1q1WTiM2dBNgDjAJCCE5qonh5+UTNZMdFRHCAEJZT9kg9PQtJvCCFu4iQrGRnnX0x9OcZQUh
hjMWeY0WzUIkYNM/a03CSjNtq/asxH3vVgGz/gzUdSyS8npdkzqdYFU/DBkg6mxJP8ITAKYZceYg
dta/6lZ/FsjqeQ4asCIVQ5aiVangScX6yjjSRDRHDp9+nASTjgGQeEVYEekogtiJTbPMbtTVrxsR
Y5PHfDDtef1Gqeck+6Jr6EqfhOUCdQHWd5pwZptT5iA9NY6t8D342XuRau07gNSz1q890Elj//wH
IUQeOXgcGQvJbtFUM4s4ONU/YDW76fMbuWJ+oOQvZWPJOXxeu97FLhCyQD9pbst4Yl/RVAWZG+Ef
SHsDtN+M4uXdylVTbIYz42JnNg+sFAhZLZ/ErifZbldbA5nZgWVrdgt5wvegRSNJyrTBTRfBGnXy
bUxBZbuDshtjZzL2coIk92SUaQW14mdX2bShUveZHVcqD5+A4Y8sgf96cBs0Yc+b9siJyY5+oyGJ
QY4CQxgqwOuvyH8NNElH70W6zo/aL3OMN7+WqCsXQqKBOr8AUYvfLu1ENnYmslQSyLB1Aknk6eIu
S4UyP25dHpaUEdQslEs/FrtCTyEONc/aKXHf/QfzinHF3zIxmrQTtO6ddQDlk6w6PYORoCqO271T
gO/QHLsc+sgBzGilsVqgTdlzu+tdTsuTPyv0pF0apXxwSZkzrPIv8p0vVL7OC0TpL1IrtWVaWaDA
7TmsLca+FuG0Qcn7IgzqTYwPTNz0n/yLCLmCe51hH2SaTpTf24JJs3pLE5VI5nZnUcnqzcRo9aSY
RQM5Hb3U5tSg2irnh2snp9Jy3c6L9K0YSQ20tVom9k4sXqKo1EXY79ANpiBWJyWOElsq+iHAG6re
lDVnkAALBMLbPYkwOLMAyTkgkah9U4tm63+JzZljsTGf90VrFvSN/dvHqmf9eeQWKSIb2WFTSfD6
5D3CzonM+9sOAgg+I8KtsOLj9wilqwgsCwiyDdPCku4AlZoStKCM5U+QAriKuhrDWXmsZWLm+tC0
/SGnl4waolXK6JNB0UzPyGOlJIXMd3pJe89/uk+huIkGTVkjB2TIUvvlN2WcyiVq9LhvZbhVs+JZ
lPJR/xcYzex9wg2BN1kaT7S6jUC71sT/bw24O1dr46SBjENIi7aUGiUN/OEqUJX6h1Yag5nJNBxN
E1+1SkA5HCxKke/QbyyvQsqYYrkZ6ptw2SljUl850OTK//KsP6dJX1ma97un3KDDph5zLiu5nwJ2
95izpzg3UR+fL5+hJ/y1DypziYy0n32nSxJSH0SJMg8ngcFT1rvlVrQudJP7eJfjH58F91IWmGxq
9Hc87qgZc7au3qTmhkiqH/gh3zXlWgapoN2Ip9IUe6ZlfzyyZ/ATB7RCXljqb6esAeF6jjlPN57y
xhZnvzrknCMfUZILFdoB54GSfCSgZqKcDy+CxXQLbXjM9LbT9kI7Iuq2taD6ahPqCek6qhq63hp9
iXSzspwedV0qwy0n+yroye2i8FppzU3/V+egFNBxH0PjSD0J/3Q5hKuogkCRMQABUYdn3hi8ETOC
Z3oTem+PWHhqx4hpflxhLRU9aPkaMFuNxaU8qUQpcWX+mas+myOoICy3szzV2Lat5Db7F9Xn3Tz2
gJFXH0bbwQZzDDDiA2TXhQvetrkfDwzHChFOqqsX0wB8nUQk1QGeAsMwpPMVfjseP2zviCICJipH
LulpWXklDrguJzwEXPX+IfN9lflGTBehymPv0i9gzp3I34UldC81tpxH4O65Qf6qH6mDVRsaJiBx
s/pm1LIdXwrws9kWhJCirLkX2YZmmf2Ve5zJIE0/OW35FeDxleXG27NllJI440XV9m0fQNO9ULKy
4rexS31nJZ/GBOE9b9DV/96JK06bLM+IaYipSSxuRq23yVpUQIFbSwkDFF6VPo63i2ql2jfnS3Sg
SQIKzJNtf32MV59OqZcCHDzp68G1cepIv3cXUqqidYOeb2ISdGToVqDltnGhVYgU3T5382el84Oq
JxCYDJ4hTIqM+qRzTzlklSLD3RVAvFhLWqKrmerXcgvm0CMBPA2BC7uM69tQwYfm0AQCzKc/I9MQ
LE28tDkQoipMlOEmXNVncRsTLZMTw9FoI4Xggv+M7QFs2nN4eTSLwKBZxTUNuX9Tw3tbLPBqOTVU
Jjxio74uSR9QJcIGClGUd5L1M5FtgyKvUPMEkBDdyzggd7obd4TFoDdPvvJ5buBfrap1i9C5GYzW
bxRg7A9etFKIxsK9I8Xuwj1U2B+Wm0HucSIGWvt5nBMGMH7PSVCnXJkmfuhOu9xr4oiWY+qD0Hqq
JVKlEIOiENke4kH6fjd4HT9yuU4Og3uSAaHwNVDIJduUgNGWYmUoXwI+eawRin9nuMGyMnikaEo6
pQJeJRqPEwRqiM/f3k3DX36CwrHFdsgwOMD+Auwyz3TmMc6BTAf+1bAYIx5Td0hcggMi1tchGFqn
rG2Mvn7nN6z0P3PQQg9/jv+DSxbo/AO8iAaH9CoY/PN0ntGOjZ2N7E4Rl8/5ej9c4Al/vi3/iEYK
vMXEniBcLUVG5P8lusOSgZ7d9+T/J/tHbY52OJPp3lRcRo2w/sak9v6Apg8MYAAd7jOtcjFYyYow
96ThEqOwWMFUhe+8ZKIfIIe99iXk/fSr5eIFgKT3VTDBb22pX+mkV9isumpKOD5aEqA36U2I+YY+
XVuCm+PoaPCMCDzvhBLt3Jj5WAyi1R0wRbLJw3o4UaoUJGbjBdUjdka3M/YvLOUn7mZuh96xnXzj
tpNYFN+uIqAE0UkbynHeGueKkceCchE54BgQB7VHPkNE8W+vfab6mYe3un/hg8FF0E9EwCHyVjvO
YDEAMb4twRnkpgqlaiDer6ZBV71KLhOvdqvr+KgkfAsMXuBSeaP17LC7GGPSpeYY2+47D/NIlXRc
YltRvPulmnlz1haGumZWeT6eHviwUollA/otyLRxys8/HbMKtKxJ24JM6wobhhI/XgrhPBaCoNtR
Lv2TIcfKwRMiumwwG0takk8Tv/9VyM5I9iPAoH+Q0w1h3K+50rLXymq/xev94VhfiVn0Zaiv9ga+
vi9z6eSbhHgnZSWUavV6I40pmyTVbFNiUF/hXLzPXfQx3hxuiVb8eCfxnV0qb/KlS5ATKrTJnIQ9
S3EJVWe8N5038/PYf6w1CeDM9s7b+lwz3TnvXwQeL2GiUN1YAvvq/p0R10SypyumCINdpACKrrkx
z3xfbs2N5u7c8MF3k4C1+cP4mLx08MON3HjL6Zv1QeRLAG1FEPdLFku257LippEEj8deR64XAqgg
voGtx9kCmPfAkqJLiT3DwZ13uPVDYvGxbMoql35nmVBFlsqUnLgGzyArzZnzbsSVtXQPn/8rxgKW
YAaXZqDk9HzMw3ASu57cemOoi481JNz6xhbuwZCuDf7L/UreFM4FI9B3mIDRiUklNrFecb+3j2Sx
VbfbGc4ABnRxbwKOrB+X3PbAB/7W469h6NOVoWjE3eRiXsjvW6IIp3FsoudM7kVXOOg5NvDW8n14
U1hIkvUZs4XhUxPx/sa2cJaRoiDaz6x2AvgsLQjQe2dJ5lwwd7CzDSNc8GVNL/Xzz8wyVogBXHCx
t5UZ1O9xVbgv5V8eKvJLRSp03WniAIz/mBXPEZXbXR4zTp5ez6AWq0bIE955LZUky2wZ4bD5LMdj
Tr2fIcNlUxoGVg9B29XyAEkg2ELExTDU8XYr/Nkybn+UQ6rl5evQ17Ha0fFVw6dyLDcHbWzwOpDe
v3tiX3OH6DeHFhHiIggjY6+gYCl9rNX4FiWrAvBSxh3a38kMmn2pDyGdhlLv1xz/ASbUTMw4l2ds
cGmUJ58vTcWpPrWevoSCNMeqN+sNrCjhIrJIG8Sb92Aq204MKwmXCSkzTuTK6SUe3ND7cMv/boyr
kl1qgEhiIkY16+IwcbT6EWe+iefGDStB2W05Fs2ff0+cn98bhAE4rIxdJ+BVkArjJjf+bsrd7Yx4
2+3nv6BtLz8UBMBXbRQjIuZuz0nh1B2XqsJ+xgcoZMCkP2zCqHbszLoSkeDDas4CHdNuWbeJ5yaL
kUDUJTNl6RpnsqUMie4tioURENEOO8EBgYuCyIi1RLIPd4D4BUfc5DCCUoDC+pWx04+sYSB5FW96
yBg0np40QFZHPvQdIFxM43iT0TeFRhjmyVpfdUXDPsvyu3zWG+MCjjl9TWxdiBu1Ci6RjPb8rfHN
nCQ2PT6ylrrNRxHQtk+kHbZTDaNd/21A/HjAS8Z4qc2/E7/QZDf8DjztfxGdfXfinQJQD0VqYlWi
j61IffHmLgV0CUbsa2KiT/uMo9PKJbaIwb/tp1KjZ7ybLji7PabaYPMK6wW61b1UHUftE2lc2Yh1
8rXGbkTrk1eWLmo/c+FUwQVLPXeVmQVNvCvVim+nxavIwOrlXGVoRZVpw8NS3LVQ8v1ySmGyJWKR
Tw3SBv4LYsxcRnTbkFuX0kTZlRoT6zCNQ8cqNbpEepvjr00QKZieGZQh/n46FeD6nofoYC7Zson3
jP6kUROTSgEGTxO/CO3jc8Wq9MqBwtlo43vmbIflAGqbehULcC0UXb6Krf6LlRt5HI7Exmi/7Wfw
XiC1PWMyr9Lne841PefyhiNLrP6fE1PhHhiZd29CaTx41vOvqWiMfgrk60p8qGvBMRhbD9rSVtaG
OnPDODCvJhBBvuUPmcx2JyicLWzegJlhdh8inEZ9mvq4FC4afiX4EM0K7iAFtLHzhSxuCmwEeniE
wC1Ko2sebOeGH89EtNsYYwQIyrhCBsHt4Z5kkOaxnBZN/XPpSUacasw5brzVt/3aluzQ7B+xxaR/
oHlCI9LYGwy+zRTrD1x8rlLCPGWWPtBbpZGdc0BuG5juyIqRoLuyJcWo3my6eGFzdwDYkoLH3u7k
bvgF4QyNRXpfUZvY5eQFkq5rqCGz4+eOs3sxx3cMP7tqxi1JEfwgjQdP/RT7MPRxRhrp2Yd4Ya3I
ev4HSp43DJSKmYs9r+K0Y/PQsBrO7JYaqX6vpkSR2sUW08ywujq+yisg2NBxfJYg/RTNWaE2pjax
WgnpWZyWwOLW86wOQUnxSY8QHsrSwmd5aEwK+je1CQG/yzeURQQosMKH6Nq4ylqUrlsbK3SH4ins
a+knHFyXi8eeh4Y1SRp4s8+K33hcWWYD+L8aahHJBgrYieoijviqv4xOrHdfsMucPj3jxIzZ3gNO
U/KG9lnviQ9mi1rLrFDU0KvBcANX6Cxr+tJaUMETQj1Y4EcvLZxZp1AYkCHiKRvUn+I6zsudu4fO
FXW2+iyWYTO+OL/OyN3TOTR6gQ5ZeH26vx8x7YMZpfH4O+VA+QaUgaTsW1WKcRU3m6CfiGgDeqv9
QZ8jZ7DHo2DWHO1rgIiDJLkC34d//43up6vkND9aqDiKL8yld5zMpkwseBLyDCBn+UE9ZJjGC5ZH
0E+91vqgIj8hgaIvm9cC+H6mQzZ7i+7sh5vEpv1zAZHCzEabuqYeCHGx1jj2c0ZFQhqMPOGCI5ya
Iyr/lAnrXbvJ5zPf2Bm64J+DG00zabhid88ZUnWK8KRQPkMs7CgKNC0+TMQHuaVFqMGxqyCLIt/u
+XvlPHL90a97b2dQKwb3CCtW66sW6D+XlAIfiQG+kK37A8tB3lVYDhy8NP/goI9OQPX0Yt+HpZaq
gC3EI0286ZvhTkVKvkCoBqdF/Nn+YoOTRmhZHEwJS84H+AzrX4vZU48KuEgzYh0xL+tIYzYNe6PH
n53jMMdB2eE+t/Xpm53sXIRsHbAlPnT2rHn2lZPhD19WHsIhzZRiBNnLsZWg8lwJcHpKLzqZjez4
L1MIROdHP8kGjoILAWEgo2eEMr2GFfmmg0YJPntWGby749nuDdAw+x2qqoLtXQVnhXM0bC7GBCD6
RQViZNMOkj4ognGyuSlqVMUr2dtixTT3oaA3JeFpdHaoSAOJJ9iFORp2WISP0PJl62XMfk9bb7Mi
oFnGuBrsAz2RXlI+VgOVnhAPlDaELXVYqX+Y/q+cqqTNlJRTvssDM5cjfXXv17QC44vWDDNKJvEQ
t9R1vFcupz7JlFJGmAIYi08jy+HTDtGWXcJdiM67gr+Paj05S/aaPu92hxi5sbx9T7DTCFwGciiw
AliNU14fDn9G+0kWTpREo1I5jlrfxYKpjB4Cga4Z59xxhnj4S42h5EmbhIyvyuI4BnxflifT5Eal
s5unvhq8sHHwIG4JXAwDmuux+e52xf2oiFglZEkZHWR1oDOGQw1SfUn01MsfjpohV3djrqc2i84s
q8AFuTu5C8FC/092t5ImUyXrh5Xi8mX6iDYf0mSk4hewZDOMCb7lwz4x8pwgZWeHeMo4BIZsrbF/
I5qVi2+ZYhvcwh5vJSaE8vKOdWL4/V2iAgykbx3kxNjLgBHFVl3Bwa5ZOGfmYfA47bishnUY0HWg
GRmL5i0O5iPoW1fzslWaClpmaiRUuOBmEECwKrL53JZ4l1CQZqyCAqM+Weqfs2z5UhhZYDE77vI2
ZoVFs4wL3c8Q1soqWHiK4yoaflhRgt5/tu7TTgx1DAHTRD2jQ5MGFODd7X65ok6GOfDa2oI8j3GZ
4LFM4+3F/ko6JPWBPOgntgR6IK9rE0k2mePYBJPTnURkw4YcsezgYBQZp0c1mOKi5/3dRYfpmmlH
4RClIaik+/uyhwbxUP1oo3CUe6CuhZYihjeAHLWo8nD+/Sqoo/DVtpudY954n1yDjy0qGyvGwsP6
eympnKdSDsnX49eaDuovK2Zv35z6X8ZtdgvUtCENYOB+NVJBkEYaNbAMzwrpef+NrBK4fPkKom0z
17Qhku4Cb4yzS/ioT2+AC/8AfNHk6WK8lPyeQQU1ToMc/qrAz8fmOPDGqwR28SHmm8QtW7/0CEaB
YMXGK6ZZJQb4k7rzh0VFSUXmmvLjP9mzv5f7CZzceiuLRE8BHAP1AyD4e4e5KRxbRkHC02NQQF5p
mNwqWD2c3QL4tWlMPatum02MXAQQoyhCrKy0awgnbKWb/1b0rIK88E8zTaUZqP5WNyLxYYgnnUZf
OQJ+aX8ri5rEHrCalcRJn/RU1JG0xOIFhbeN/wqjjQgmPSg6IlS5PMON2qlHKb9DxDXAemzaN+WX
6GMoUzM09tj/BBfirW0XHxvRjU4rtPgJFDs/L/yQJ3AfuKNQERE0qISg7iIAb1lLnpaFSYslkNFE
oB99CZVUOrzxCSKsqaPJQJIs/AF+V7OdIyBdQdDtkMZYr8do3HEelUHbVsP+t1EOvKTeZcBUosaN
nx3P1tbJOZ9Io8WOVSOAiGMLaBeVAqKtV+PPIEyuq/s133hplfRArHcamaBCgvsCHKmGqABB+p2K
yXS8TNggfvxh6XLPeOhXwNe4oM6I34Bx+pUMp3+gQad8coRZx05WKxUTZSLsOhkgJsQoCRF5LZHH
+G3uCbPnHZA+AkPoFNJdJULnqWTW/ePqfQTgPVPGzwzJleP0aj1XIiIB1CbsRg17bHqrC7CM9rAo
Yrtc+BcQKL9KCK6P76VK6261yo5sLteKDdlDa8vdJ0ZQRG3kXLSwv8JHTkD176xB6nApG9DuYqCN
45CrrHnJFmVQ5yaEHfSYTaNK9rBzEqtmvYbhmFzKDB41WOF0sBIiZAZUmK3J+xPV5Jd3AVLz+h7M
s2EJHZ/ksCo+fw0Vd5/LoJKdzGr9KSvFdG2xQpzfjmvpg/JBsj4C407SEposW/ndJiGcynl6+C1h
av1AS22qwQyLDyLBTnvAcfU+8+UZypiFKY0QEPbyXJ6nXn7w0ele3f4Qqegkg4BBQIpm7dcBkA67
rvq7X9r+kvpVJLqb5UW8Dxq7KKOY8LH+xfhx9ynmo9RhA4Y+rpr/QhwgitKHKJZXXqNMaDGeV5cR
PBPc/jm/9k9MkGQC2ogbJk00e8W7qqOFepKG2Gd2fmKUl1WUrpyDMQ0F0aB6jmbIDz+6IRrLyD51
JTMHwY5ULYZgQm0CF4N3bzHcal26zA8BQd4f8CJfBL5m8BuA6uQWw5DWnAARbsIMvnyfe30fFTS8
PNSxAlzy/Fcn2n9jxp3FRll3EYy2iwgi4a1Z0zxIHXOTSqiXgXKYQHfkbya0XcT/eNBcon8og8AE
unxVouQyKW5TKi1H50Ovi0EEBxgd25kQ1yyb1zTWi6NZNFCO8DruIwHXJzZiIsT67OJgm3W5YQvh
AtTavSF2408bVxUgZpf5kqpd3JvpUI/5tWkLsHJd2ga6lX/LEsvwDpmEii4T+m114uvU8Mkq79kE
o/Efb5m+2VBJ3qGSTUT+TfueH0aKy0DPtH7W/AuL2BREYohljNu22E0MtBTn38dO27LD1N4olwrT
viuZpUggaYrXE4q5pleywOB79Vuo252CT+dQSHHDJeKhO3vUSadgfsPMmfzZZai3MFlWU5ub4bcZ
K/K3Wrd/lZN7GZt8G/5NaJtq4fdOMGUJnxQALEkqP92N8eWR6S1Sm3bDxsw0jSVzmDyEzAwm431l
po4wKrx+UlEsa4N7QIVVE4x0On/BxqjV6UMx7CnpYaAmNsl6IdbutgahcbSrgQ3JpCmOTFrMUE9s
0ZeF2AVNoO3MC5VZlpjL7/6SO/Lc4jtvg7pDzZEJPJ6DvJF37ePuWTzDQxjZb4wtQPqkQdCvHS5j
mGV1q6OC1OVDOzuxwan2P8fG2mcVIx6yewJuonlchLJrjAyYG9drnEJEmeP5Vu0Z8MJdiqLOHq32
/Lzp0/kvZyIVdcpylRqNBTMaMyf9PTY77q21k8idY9UA1bchchmjD+yDbIyWpVfk6Q07jGoL2NYc
rqiV3smDk4bxB6IXsdT1FlrkmJwkA4fDj4Vq3ML4A6tl5HbgbeQppF2DSBBJQ3AqNRd4keFHqlTl
gbOb26tcjtf4LxMfUf6j2URkHxQX0KeRUe0MvwGTXdpT1DsHcv05pzKpPoHpmcbaZb6jzzv4wsX2
nVZcQ97gHfVZVPU7OBDS/zfH0hab1eG6QxpDqjREzrNilc2wuKJ3ucbh+NHM7KCPsiItSXK6z/v6
8TZNlkGBLeaEfufwjBWveXo5ZFyRlljyBh24mwBR/t5hfQwt3CeHc6tg6IIUho82b1JD2bkac/qS
7rvfB05iHrVOrU5K1RzZYpx/04rYi7VHzp70IApuxPzi88mm3W+2NfaKJdLAtCo+rqGmXHC2AtPk
YXyD47C36FeBooO5P7GYVKaz1mnJDWfdFlSeKzrnb2mBSkFWQRDeYwxBW7IiDpM6SjMCl8ddFTXf
XV0MZCfynjzeJugdPGHolJXzdeZs8e3v/hKGPOVTPgOXCmXyTJlbG6sjG7MTXCfRjw9aFHl4Hn4T
1cNt1ro5s3VLVUihAUbWouM4w4e/SBQBEaaRlxAISgbkZbfXGC0M+xsaspAXJhHtt+0eSNCffYgS
P24fVh5zGbEixpO1uNoPACek8B32kjtm+BJRQnOQ01wxSJHg9y2ufXHTFxxQnMYZw5T5dQSoxUIC
xZPqSqT6dCcXcEc1RyIDcPDFMkATvnrxQoFtD0ftOQHBs0th2WAwbWKuNfNUWlB4LRHgCtv8+DPb
6oRqcYOGcfgCSEiUe1J7Apsb0Y0UcDilkqM9zncz5VxVVL4GoztqJuYJ2s6C/CHXMhRssxNR8p8M
MxHGVdsunwMbCHXvC3+tbKip6vafC358BgRUv1BPY2ASapMQBL5+uuXr9OmyJZ7bxz1QfNhMyV9E
aowHguqDboKMGX7hNX+X+ytiJhJfsenAk+soOZtnVdi/8PCo7GVRdTe1uosYQf/fRUPOQln9Q7UL
ebjWTrwV91963eYWLCon+XgMjbUIeDAUk3oGgC1ddbEzRXAVNo2L8B7yZWkPXVL5+PNORZdbPsm0
OsMP023qIE6o0tn0dIOoDx1OSrr/G8RBBax8tHYQfzE15AbR/Dc0IgAfpmZMzN5sejCezvSQWQ7j
x5DvC8faMRycTtqIB9zhGexgG+sKCShxTU0VDYyqiRq0liSuyxrjiWTt98ZjgEyoOS/d3m5FT0l5
VYb7RJYdIIk+W4/FbeiystK26mSP++18GipZsMVmTV/dcGhhorz7DPrs9MXyI6gNE0vWeLj7wcU1
5zNDt1S4ZgnrJcalc4Ig25HHexNGD0BPb9GwmuZ0zUgfQtRzyXRJdo5X0YL5pPOeThyNsxFD+ioQ
x5LNDFMcotXhKZCxVxt2FZUZEkvmIeVCsIGDxqbT1KpXjTGWWmGVEvZ49l3l/Z36Q/MXKgzferYg
yJ+V6V+cPuulyKfz64g1SF/UYsaiOCw4rroNy68eStf0DVAIrGRsRZQHK/njbANj+lnF5unxuHgm
5yU/EtUtx/8PHtKkugG3YwXsFVqNW/BXTI7ZsBH31dAvu+A+OgKu6CDTVYvy+0G+jrZXTcZ8QQ/8
wKLAkz/PRZOz372BEAKAd3Es8wU9mJNeWTvd2b+FY+5XzVMlIaooilu3ZqEza/5OhnoyNgZ1KstS
4C77Ll3bUQ0mnmpV+AHj5RyhDZ0FCtNsYYRzkvCUIQPrjaHED0nprwxWzUFS/s2m1Ap7xeNEyFqN
LI6e7CqZcBj0N/Q5mFlJMQGZrBtqNy9Rd2dsYx5YA+ewbrasRd7SowiAjF5qFBUEhjao12N7FpUu
EdU/V8Rba2KBx31nAp4ollLwPT0xMe17KEMEhWz9Yx9h1A9MTivMvc8n0NvJa2vA9d13wUhpxXzU
Z6BEfXM1JEVhoAFipVcCoTmr+wqckONVpK+kIujavnOy0CzJyREsi3JFWg6AzkUbQmKvzR/obhox
u6LjrYmo61VB98HzSD7wJq3Wd3Cy4Wtc7SLzFw9mke8sY+6+njZF/4NNb682dTI6LRtDdAd0As21
bW6/A1XUvMBQ8C23BwADnYHkFwDrjJCU7vf8rNsw6nSQiUSMYN4dVf+uI+SUJHikEUw8J4QBkvET
xes2KzDBwXDxOS8WJ3m7SD8Fg9LiW95b3WCGmfP2QQAGUTc3uEw+c2CpS+2oa5ZOBfzkjf1ttJoY
jbEWrWkqJbpxFdEZO+LkNt/ywtQFdx4gPAmbv56bQ8OG6yMpHUwACk+ajxLZatykfq6XexMlU2v2
6p3i4GUBAnPeWxT2/hqn+aP9C+50tJOXih/VErDMKMgDR0oDpUqodI6Q3CpHJbIUdvn7LE2zGLAs
PzxTxNASrm5n3K0ikmgskbbp380ya8XsPQs1lxiuICBJ7KpYGbiXwun0kn1W+TlIy2qUc7+AEvPK
j3ncoQaThY4RAKFRUfGU9JvvrB2TWRU0sSVgoPXQJDr+y2rDRnFoGIKmhdywSuwFbIyrX5yQnrdl
3FN13JHp/DT9NwlEjR2/Vh5NyQj43UF/jaCEzfmmV+F4aXsFMAcuDwak129utgTuE85ngZKIS56j
oZ7ETC8TF4d5hrGhEuyiDI/yJcjxJTzoFrla15pCQhcABO6jdOBjhAlownmlkJfdO/QVDCt8AstF
9blPpk8H+/3R5wrWZF4+FdkiaVrj8wwlgxJkGVuC6jJaCh8mHlhAcnJhjgPrLOR86wDXKtxwtiMj
aAUcLYM/OLQVhcozEs5qWRr1OrbMA0VGHleRe1bbY4f0wDL7ke2aAhSqUlLo5lWQA3ymWVtPA9tk
R0fj7v2M+Vr9Pvmkrs9Y30JYOglHCqvgMYxPMDrjKlJ+574/mHHXU8C93DvGcFoREi3k3wFMkdiq
0P/bJNW1Uk4wYcR5BAhHvveSlJCNBSuRV/jV5yynNImBk6PyY99aIgLqoYa7r4dnlP9VE0PmeMfk
d7aSaXSE42ioXMK9GXgNR8wwjjt4Moh9i1ukpHVf5nx1NJ06f3EcnSdliuq73JXQLoz4myWt869u
cMT/B1SXB6DJqWxcXE1/y5Irsl6ATvA8T15vlP3Zf3bZXPzN52+CQtGRn412AsNhAmkV44DKzcC4
JyeFy3Z841ngQjIjZyPy1gDwTm2zCWuzKiAujS10idzHclnuUWI8D11Xc3uKN6APv/BP0oEIqzmI
2SknVG4zyFKI2MOAplkxCM8BUXYtUth/3B+9Nv0rhGMSQHKzZ8PJIRLbA/2LBF7Cl2NKoFxr2v5B
cI2956rnQl11am5isE5LBLSg/91hU2RqEOo+90Fx2AjQCLqrZRScqN7JZNCp82KyM8E6a/Qd1UQ5
efVQvoDQ/ULouaoL+a2frX6Z6BYxBNjnrv91kucqfGY5jn5Q2hwDa3rBs1lpsomRIp1AoBGu8hSA
B+eezX56FtPuNu4LJsVyMM+kOTn8ZN4FKInXoyUoQ0/XPNKPN9+2l5H/gm+c6FMcLYIqnvbepwhk
JwnKWrvbZmUZNRl2DzRe/OLyXZS/7bJjYXfQoCgXnD7hAT7jsNHl6Ep0ABlelmn4Dm56MvDb7w2j
73SVtbt00Bt4yQDL5y69tq7tF4lCApcTsqpQ6YjPbS7m5nYjZQT3iuAL8vlB2RQ4fe8fdhLPfTQL
G1XJzlmMlWd/xCd0LGpvBhxv4SKDqrFNhEq+p1Hu7+d0cB29eIT+LxKZ/yCJcs/R9IpGaWPQiI8F
9eKzGW7FxWJR/AxFQf5CWuybuBzxGGMdAitBvxabB3mkgqgGF8rC6JyVguz6JljqtsqmoirTqP31
FoyKobYzMO/Zbpcu9OlNsicpS+02l5R+YdhCs3fUwckno3CTqYZvv7LSxb1ZTT+juZS5N6zlEOMk
D/BErD0L9vvJmm//Y/j9CyLdJcEjX5fERxUoxMo9cjupNF9X9WQKnlGcaQbSFTbRpS5ZCbBD5+SF
K4BadE3I/3n8yTvC3LKuLpbn97/0MOYNYjBDvpqpnykMQxUK3nEW4oPnW4957M+XFSmlX2quraxa
gGEG3PEYj/qZb5p/EaH0l0OJonjspYLmi0RINgxQJMK873L/5P2eOsmcFfmS5ZS5no7tiFP5NfEZ
7Kys6SIplQ9kYB9MZGBaX2mUgnpRjEzMujOGrePJST8BclSaibsZID+cBBBELMHvRsFjM0Mjq3nA
YCzZYrrfIXMAOgqDB3paHIMYUF0RW4we0docEnzyYveKlNZG/MDONeu+MhFkpYh0rTCoizIRlaX/
wO61fLjk9S4jng0W2pwYdw39JXOAc43fz9824WuD34t+e99uSOEwxtKIm7EHUha1e+JfuSjvzsGc
6DRGNNqIdSkd7PIxIZdeIhXCixCN0VEiypvNoFsik60QeDKSNwsnC40zD233gm9FGfX1QCWJX0FZ
PyPi77Y1aHpgCLhNFRypKMFfb+Qv73Iln8reh0xm3UJ0Lquxmk6nx37JhbFZEs519X7xTUSvCG8o
Ea8apcUy14/+aXldw/EVnogCbVAAaL8pwEHkclRu/gMdfL3alYBZQjmBTK//PEZPW1T6nMTQmm0f
BsheK4zLJvi4JaoyF4osMpWq8NnXQKWxa6Fcb/3eaMVtn97q/7LXXH5CTmiSehO4dfeDLCCrnAcI
T+qFmPlhivdm0Nfa6Pz6UX1GvwIPz6MLMfe54Sj6YCjj+PP+nvQMEGFz3mJH9DeLWGsfMAPvhOOj
lMb+N+71fIQTmGZnlKjZq3gswHECrRhVb5z4NPgQLDPyY8r3iD90hqKJmZZKR8lsqLw71G3reCXu
dv0ZmSXCNACF+s9Cie+PjdWgSZVBEEEexC5w1IU+lsReXRVDOF23qaLT4zuPWTOHeEZ7/niFn00R
BUligwgz8WBTsCYYTyOL8BZA0K+FJBoSdhUJRKXhGU4KHk4lVK5sXYIEh4W/5MuTT+kzQRfPJ24C
zOVpbkqUsTSel+MDzUEgFK+rto9JkawAd4tiMiFVmkmc0GA2IFLKuACnViz+s3nG9xFjidifGHsy
Sw1CE10+TPXHAeAIrPCi3FPPVqJOzuGlBkomlBoYAmHanPYUvDim7Mvb8T2fzVR/SFZ8qCStMgKE
uskZjCrfSloCZ70PMZ3qL1ohDTuVbywJ5jkxhAWBfMVmK6N+Zk0cZeuwVzdf9maRoPXCrUt9eDPZ
KFlZm/J0cZOoTPxvsvQTXYpJaS4AH1Rl4qXnojczX6woKEoVBXxlEnPQMjTdOI27/YgYr38dzRUR
O6YzkknSGQscQ4NcrTvdmVhuTeJ8xo/JcdwfXCeUbTxfnakf/S8kSbXEiLn88844o59e+UCllQ8H
rKGId+wGCQvxylspTqhAs726b22oLQ3tRWXI06vBZOwTXQWQcQuCBqDxnooEav/NPaiDsODL852D
bGFs171o111J44mZXdAStda5tgWtifluvFhkDUtMN3DlA3LgyX+3wFevV4+p1QcjeFBPN3Yq1Pkr
CpZYHsaGbZIYyC3vNP1whgGBJeqZCY54TGTFbv18nnhhSdc5sc6gYEzKsLqCgQwqR8qHICgzIllb
bpf1SZFjOmdF91CoXvALar0U5TgPOZr2I2ysRRT4fbUkIurUlAramyechNGzqd3lIsVqgbfkWq0g
Uc0pZja/go61a2vtB5/g30jQJ3z7jCrrW/0pDFNL+tvvDCCTPlL1q1DMEbbmpseqFS4perLPNxqn
dUvyifH5GSr7191MORHeMOCDH9dBbRocrmMgVZOecYl2TU8aQpRRjf8xB5RLvifNl2nWFBMWNEpf
TZraAmq7sD5DOHZ4ReuwwRA8DiXt2Ak0x+apjA1K5e4lsFySZeqh0ieyyDt3qhsE6HGyy+EgeK3D
31XOLWEQF3KKm0ekANjG5QMqfYHgUCm/iRhfaWOqmUS8e9rkZOyg2fN1W3ZPJby3dR4xS6O9VLP0
KG23515zfFscWVVmrWLMkBzamLxYF2/R4WXYkU90cbQfy2YRxycQuJgpvi/R2A81+tN7ZuxG8Nyh
2cLdd2SFHCU/E4d70p6onVBnvOpqQhKt4dirZyKCBwqoW3cgm13HF6l7FddzE7sHGDyRxgIvKb2q
I/AfaEyG5te/2LsAegke1bixoLEx/wTkWdZhow3+PyaQYok6RvnFhkzp4AzbYHF20cSNx2c8ehaT
c6XPz9rtexPwMc5HY9t5saW6zimPoG+bIzVlqUbm1kHaDHtOc6LZnktvqsNLP4R6A3T4Wjr8irfm
Hvmf7azGAN/bemJZvsiq0XlDJAPVcx3P8hDmprXxFHtYYbrDiGkIPx8TMsWg4DIMtQ5isZW1ovM6
3dALTvCY5tzGWXzrHg4ZS2qffuGuGN4LD8MQAFJVRqlXu/9ytDTFOb1Jl3OgpT/3imjXIFuj5bna
fW0kDwfrvXDNSya4FpAQRNnIP6ki/Ofwr7NMCuCfYcmPLQzOlW48CP6swIoCvMLKU9/njv3wjYaq
LaEkz6ayP1SuU03zrhov35ZWuUuBWyPqlCj7yC2Kq8yn99Z65ssohCxtnEfV8akimJV51dY/9lMH
RPm+Zf6oCBUcY4b+kzHWXJb8z2PmI1q/kQdHudksCNU7L/MkKMqoAuu/ZQOcPEpS6UrQlL/6UVAL
u3Bx5jDHE7t2UjL97AjmUHVz5AITQa+dyQm4KkH38ejhfg/RqXhqzJACPeNtRWl2G3AR2yR1tMqB
QBCd/+2eBr/Ah6P1yrFcfmBfDTOoJNun9KsuKo6ohK6x2VUCbmOz2u3MX5jA9dyIjd6IoWW3gQob
Kui+Klh2kvUs4JRkD1d7AQvDbr5Vc42WLSaCEBjbee6g3Wzqs2/Dst0Eh1jTwWd5pKNBQBSJDQ8n
Fd3U+gkf9iQWITZ3h6tyfRm4H17Y747dU6aTlqIpzxKtxkDqW1OyxduBYuVBd9qjbVVpA8pzah1W
ctrCC4AEVIsP5XMnQ9RUa68zsRSShRep/cChwLQCaRyKNrt9u5Y87zPvk8tLI90YLxN+GfXuthto
UnqMgtrYV8Q3PWGEpli1O/b+wABc2HIJfN52Xntu+13NTgCYuowUOS2WkO/Ah0YoBN1FDDVW5Ocl
oOENNnY27TZt3Co8nHlfLYjtmzidjalbr3AxzX0Lr83P1xjS6/vH7dC9Vd5IGKOkNgIqwlPQwhAx
raX+Z/KJcZuI7qQ+k81yAd0NG9ZB61XrOEwB3vlT/RqdUaMwxQ9uJNnuCMw+3G/044LY55SdbINy
k8N2ETjhh6bj/onjsnJVvWcz76w9CLy0QJU9pJCT76Xs9eQs/76Z59Tjv1jgJCkmhJHAFjQg8trO
6oCM6D7MwlkHhUorxGCRAXTKFvNITvF5xa4TbOlgOcGGBzwTC7o+cZqgsh0kWk8Km8SYYiHQZLx0
FvMw5FSAEoRBaUojJqhUNPlOiUHr3jDayFUOYGbj4WfBIQwPSbsW2JbJhctyJXg0qlG6/uTQoyQT
+BT7aITpjEF8+GCQyOGkd8eVed1/mgnVBjtYWZjhwbVbOAI4sRqnVgXMzVAFQdk7OCNri8Oplzsv
4LxuCUy45UDD1FG/0AkQtqa3i11TRUc+/xhj/FMeLXPQNZ+3WHc5koTxcbc84UVfH2oWrOeUXtYB
skYqh6ii8flUFEo4pJswIpNGAQO8rnjLleJclENlBAi6NE5DeUAwzKM9Lk1oreiF7BDjAYme3F4x
Hdax4yjzT6GZE2XbkhouK/gdpbnZm+SwvhxkZILKt+a4iTDCE4AFiECFWhSsIFRdRHuxsw/FjLA2
KMILNo+nNM1qII0XRhvthWcL6tN4j5G+dqEHjPoN5HeQokZTB+7wO01bwaxzQ3oHHwph7ESzKpzz
2nBPKfXhk0v8lqIaxSJz2IVifiT3ZXVYNe1ISUc3Ax9zzx96abypUpyJj6t64fXJwNnEY7N93JT7
iWu33wOFuZp78sCyJI8xhsauPPdcuN0Hzjd2XOqSXNln9MlgH374rm01OaemIrAEcSd1X0/CsCtq
JN0edPV44obva/X6M2NT0rcrFXXdP0YmIwYAkyEDgVYWaz2MxkbnJ03nrgVi6IP4W0yHZqBfH58A
bEakUrqqI14f/SeO9GgSOPbD86uI5uqqWAHNBhA8zRWPm+nuQwuSDSeu0rZajpmikWnofERTV1ma
onJU2xOv+TwEM3Yo24EdYeEYuFHgqvW6KMKP1hWe9D1mb6TciWD/OgS0VBmNBkNeRxo2b55BoldQ
wcZmyeSlmj13SKwgCoE7jeoJ24UJeGKw2RQdiiH0LXEH5L5j0WHOO5fJ+OMDYHwmKbXc3pAloyl/
406Ah4yxa3GQrUr2UhFhET0ux35HpxB3w3vBY8aYApsFJJuWTDtqQhPZy1C8zXT9clwwSykIyg4n
p9tb5cHWF2oU5jeElIY1rL8oyxW7Qskdps/43bhjWyB6BNX4mb4M+PZ7csQPLGDGQJJuaAEXIk+Z
LrK4kpm2LYIVVcLdVrhJY+DURfNtw3IKN3/gSwdPLcHuTBJzBdu1v+r8v6iVYs2LT+7ZboXR0VOR
GObaD2naqYWvIGQQQAAPrsfiBLeAAsjSP9loMVhQaXs1cE8Yia25TM01kNaidf3GSkWQVE8jhv/V
EBovF627K8WO+QLwhhBhbe154O3WmVny2GVj2f6RHmFnlqKQG5SL8ty07voN51vwUP+Fv9/WDTnF
dOBtjsgvDuS2yln3o2NVJ7InECbS6RP6AiTbYnW2+cSUgXU0FbqIeRo5DwU+9R/zxmtYSzFtMyhY
E9KiYTCr6cf6m5y20+LsHxU6AXfnXCuBQEpunu2yOn5pcMquyEOb8twbiqTUyK6xG6qI7IDdMwlR
smkuQino1x76Jp2SDuIoL0gmjjF6kW1qGv2lPw51xdqLf2AUEePkgcZX6jRc+Egv+kPxHQcD8Hyl
SlBsq3bNUCeMW4hmLRctDP7kYRH9i8DxOiVrbaZ6u3SbI5l0qVOa76T2gVIihruY10sqnkaLN/Ae
Osb7vRoi07d7+YRcc9e3qDIVuw1A2z8/jBlCOb8/M2HWIHfNR2lK+Lejsv2FfXhfoOsrBWaSzWc4
NqfGaa5vr8DjNcs7Orma8Kmf/w6Y+wZPzwzU+DS+MudsLYUgPDPl2pnDkVuFASEvHGOeMyWBFtpU
SqAujdAsY9HeTrfLYgL1+xWe7dF66wmb7xeyPWsF0k4ms/8Wd5167rgXqvy1OQCzVA6ErXzPhU2o
weHZ5tRiFeV1+Ap39Oas/eZ9fM+JQHJsaz+DM6l9KXXrZAvu8P3Mu/eJNH8Ve1MtJrcNvdQLlBkg
qkYXqTs2CP1C1ImIGiKUdcfF8iFjryUKJIOL1iUjfbQVYSwr3082AvOSoXRE/7gTTL3/8YfsxWF/
PegLg57URqpY2EVd1KfmBWvnLY2lAaAz5RAECVzODoSAZi4jNswIpuq5KfioGrAMund1zb27ok9y
gRoVpCm0vaRukqOUC2W8bSGeKaQI6c3luwqZ686z6Gl1YK2oPzK2VHHUUpchP1n/WMEZ16smB8hp
RIRW8zEOtgLkTAcuoc6ZQ4T21HJcEhGIhthO8zdjUzSBB5klxz1gd/lUVICBrlKr+Qe/uu4EB7Lm
FYhqOwqOEhaxt/611Vl6i+VONibxA3POrp8JjVngtgUeD7RNaS9x87aKdkwUqZg12gJTL8WeynzW
KqjBVvFseUqaxcGi7VICJhavpWLIm2fxmU9FAFn5E3RdBcWKK5Q6reVlItE+/u1Zt1lx4IvAf9qH
GpwfkI7OwlMbNZJRebxqLC4pVqs6MUPQA3aqYB0znHCjgIZSkFXWMSyEq2Dih8H4MJ4tEWoscLK5
ae7FPJmEYoEVBBDy5cvun0GLKE5xxrO2SseLf+qpJWUpleEtVL4s4To9E/TWq77SE0HFueL3WilA
rtZgJLTAzrT7ywvoUhUY35x+cp+nSnS//vbsodVzqlajPXzD9sug0f5GcPOokKSdY6C6GG20Sbyk
PDofJ9jT/CRWBuH/bfcqyJV9CHjsx5xsYf9LAJhErtrdMsJ06YWVvNHsu6VbAYr/ZdE7D+7EtVr9
bPU8Ciayhe/ZFPHkLsIhelAzcCO1eRt6d0SDpWU37WPislvy1wF/0/IDSxQSQ9sfcHKZnNhxoyb3
xJqgZzYDwaxbOWFfUHPxgk0/MGvcDeqZFZusEKsw5dYbKzbMb3wYVkdDRMPNEEnQLQhL6t8BA2Tk
KFgqNIibzbxyai79BTQ73i2rmESlaPWlZP0zfZ3TAXBbICGeg1J9eXM5Bln2pwM/TgnsBrtwzk5Z
CK54UlI2sIbQasxNMmv/g7gb6XgBKjcK8PtWxOvCxgth7wGg8QiTPKlk8+EEyhzQW61CKLpsdRPj
HKoIBMGWU2kgTaR8Iyuy18zBQg8A223dUMWVRFcEjnQuilXyQG1hgo8fq+WJvUjw9MVz5Cy/gRKj
s0K/G9BIfXasqb71WAF1b/MYADrKMQcgInNfKN6RC3EacQbnjIwoq8C8wfkVHCXpRGr7fIXAPLY4
6olynL96ItIQ3vrJMuCLp1Uq3UmvXBu0N3bEcv+XweMbyh8eBX7kRamPY4RcVu4lK4D2LAh5TD25
U5fyHdbTZZlr2IoEq28SmgNra16mvUdC3yBREFqBSbC9rF/Y9AlgPG9OfgvPmDPTZ/Wu6Fwp7dwT
gu5M29Hbh0HKe1aLXg79P/++D2bytAy8H/X6XIo0KsomKU6zjtA6dAtG40AF4hvQ+td8b/7PRQjg
hEZvvPgHtgDLA8g5OBVUUrI4oFCtVPhZUwacrpx7X4r39t45EkiQGMSHRhw10j0v9LwPEJ6u8yci
ckoCSn904ExmBYEHLEwtOhg5tuvDXcVUzTqqoxJftjyKtn86ENQQPi1hKgZWq8BoMS/2xBqlP+Km
k9IMYRCl6c2UNQngESHCfD4ZI4pRrDTq2AjMw7KR5ERnHcco7GpU+bNQaEAwC59jlSpmnOk1WK3q
BrJu3S6wRHXri7liLfJ3CELQVg5+0rKqXJOhGvNhRSbrAx1W8KgFcd8kcgf8htZdWu4wsBFusvGq
7g0VkzoSY3ppFHYnRD8Fjy81IUqZrz1d3O7gwK9INPy99J1dQXZPPXdCdlgyrob/ixHbWp9Y0FYz
jUqKhr71+wkZvmmA0JV90bI2G1T8Apj5Uicu6E1sxNkk31LnmuRK+XcDSmfx9Nq7G5kqdGZmGhKs
HKKp8LatQ1W1kq1CEFTwMPHG0tivmmHSRLp5Yladr5i8xXd3RhuXwAoAV9eFHIYmMI9ePrzO8I8A
adW5iF312rE1Yf6FryytIpvisk+C39Nn9JZV6oFA45QyRO8VcwmhNLRTJ+gsD6jC1Uyn583oeLPi
Xsa2YL0O/s9EMiDPffRX5iUwoL3MXCYCzLRkGZmGBPGJoLLoEwAOS/h9aU7pEpHBMfYwg6F7MP/H
LhZ9/9VQdKD85lRi15KLVYll4K5/kcqL49UObKue2pU3+NP/qOYBHrd5VJ8vZQTHABD40uAB+Njl
Pg7AJu2V8TXL5gBgT9zGVIjPLPsXXJDRVPQVKj/YxBEA+CleIlaxS2Y9MlHPHmL+bDrk2kUC4I3u
G2uJ6FUxbpD7NssR1RgtX5OsHov6PK7xvkduwWIKIVwPXCIb/u10CqpTZIZcv5BTpQ+4VBSEg2pS
2Y104IuIXKuspY09HKnAMn3ZdyH+X60Smw6Um2l7p1YwFpGyMdfN3NZhV7RZzu7nyXuCqWAZWb94
d6yi9q2Wf01Czp9a2a3UgO4kXgBmDenKJlwpQdo+3a2PfH2omyXaVOmF3/VXgNVvD6dYhZXgpSVF
9S3upSz/9jHDrNXqmaSCg7Ps/HZGMtvnHJupz424BzlmRJpD1VO7lFOAfjBIXzZmNlDpOU5/FNru
7+4T8Zqc/C4wChz4TtPnAGe91sLfTJA8BzBDkiXm1n3tDMEqK7nD8fK7O10+diI/nQJE6XeqJNid
lDd5qssAM7BSrQEuQU78FGFerhfGKqPW6dNab5VXaH4QPWzSN54x0l0WStwRX2j4flW0dRJm/gCb
V37kSiNOsMHFPi2SAGX9WWYGmcQiv7B5J/GpCAIeJ4zmTI/MbjPyxL3Bp1pDb5er0SEkrFe4izeM
uxUkebTCpQDt+e1tI8HVZ48f8VU10Yu/i6abxgMs/yVdVEd7A3fGwo9Q4VP49QgUuWx59zexiAxP
lZ7b4DmNje3qBLyMSwU8Yl03uBDOZ7ipPeTHFSeepteK3N09oxpAEmFfXwASGGuO3/htGMxaIWoy
HyEuzElOauQY5tiHEgqYzG5DqTQ/3ixpsOZUViOyAhgVRC+vTWyFeNMtYS7NS7e+R/GMHmw6zpa/
TTT/wK9/W62EA1nm/FfPkQ/7EDTTFVPOxxHZWvv8/BrPYFd/SMz74n4UMq5gRK+7vpz+YJX/k9Qh
bFHtLRKGH+paBKk/p4Z9F/BVyuPKw+h2mb46Z/sYeF8uE8pY8AzIBYPkgE5cl3h/jyJ57tpIjwp7
yTprMalYEXczqrlrWe+FW1uhFZ2r84uF8PHEqwP3kkOva8dNNuT65N+ecO7aDswQAn6CWPQlnD5z
OcY7fw5g4uqNWIdKIaixpKmArbwxdc0XdWG7jbdgs/YllN8UxYrvms8JhGkfZJbsss1E1/uw5mF/
EbIRyiY9jJV78yss+AwnqUYXyWa/9LoePgS0bFbYHQBDU41d7OV2xiMPzaQzymPpG8VZqH9bMU4Y
XT4DSJJ5A4QMqcTcS37UQp3JaduCjjKsFKKbIkBIhMDxaQNEYKNUd/rcEVp0z1QjRcx5xR+58uan
ZLuojrzef2sdHCWfSYvS44cWi05fDRpE0U+y03RLoRW6drKpRRn26n3ntK6ciJBjBmVFib4DUqTX
ChJ4WJvOY06+r51dkKBA8/ES1otG37DN1lghWgQu41FyuMGyk5G+0ye9c7cFW3lfo4cfNEQd6TtA
8kTQUqYeMkjHTOdKct42l4xlos+JQ4I+gDdjj+n/QlfzODu2D3hZzcf7Azk3DOqTr1uhDB46AQV1
CIGg1Obwg2E57nDtSk0X6lIinC2xqLSnw1YACiwH99jPF/lX5JsUxDOYJe1a8veYqeFRVzwn/sE/
cqDE7nUH3wD6peIlwlGo1tlG9aPDbwnjczsoysplNXFFBwcuWpU1BprckIVC8X421d5d/cayDnxZ
uytbgvkJmXX2U8ywne5N+6TcVS6b5Q6oIadfI8jnzRGUQiKq3G35WRFaFXjenwCqhS7MaOe9u5D1
8pTalHSaBETovyEYFMBVI3vsuL55pkFFge3m58kRX9XOhARH1stNZaKi0CE7qzyEdNtWOxESOfmz
tdan3asuMrxM4LaN/Czos+lZnRmemxuYVI9bVXk12Ss17ZHXEWo3/hiH/8Hmyq9UA1ztyqH9PZvw
Z6Uk8k7oLQylrlgApyB52t6wTNrJ7WzADhIFQ5WyBQXCRZ28OcquzdpcbzoS1NetQYjmxp9W5Get
X/UwKafqB4wRms+iVZdh0wPWmS43SmGc5gqbtedkcREMq7YHOLlqSo6f/TPo2ba2o62WKOJUE4vx
JF6/v8ZJXsPYhdJzwpaB5GXXUmMmZbSUyoGba4bcWSffrjL53UsCUtPWtsQoLCm0ggrKcq1oHH3W
nfCbD9EAlZKfLjHJvnMB+9UjfEoqs2anNTR+jBaNf1NuyAISsYJ47geavnqK9QaKvOxL0K5m71yr
IunPOfdDdqgWg1BeM6b/OoQWBs1hKAOgXQnvtDV68E2Fkk7Z5qG/CwlWc28WjCMG2SojUvqaySYo
vU5NuBiA8Ka+WD2kgj0JC/6eesvz79YGjgusoWIKgzJHX10RxRMHVCHr8fxU30C5k1mO5TGN0DWG
vVKFTeLkAYVMhaCKz0/ZyIuOn7aCymuKVZElnaL3eszcA3P9yNBkdDgdGI30e8Yese+Gjs+t+n1V
QmgBWGXR4EBPNfceH2jUrM2vNru5YtTdQijoLf+ETq+13C1MgiYnfy8dwNehhYOzIPwWRxZAJF9v
w6+nAeZY22ap5bN0rBe9XPQGC0vy5XcfUjJms9f6LPDmH8NbOAyEzvpeG8Mpyt64yO1vasydDTlz
5fz/l72OuN4hdTBlk37oesfAyNH9EZb40A8xUnN4i4LjtSlsF9mX9w/3TMIQlmV3Oa2TnjUH+EWy
kopc0ujiITvt/LJ5MngLF0bQeJeamFyrYrjSPK6VDKB+4D/wHWduUJX+lnqw7ZYOcCWwZYkfCFyc
fGtl3PgrTx2tKVvBQlxrJgEkzAMHHfPZO5IrU77pBsPCKIScINJ4GPvi2O0ljYrvjPT/kKu8GVNA
Ra2Rhh6YaUobSpuE/aQ5kPDE1fphDN/RsB3b/ChceHcuhA//PBgSSC5Ev2m/z7sI3JuKXVNBXqDt
wxzS/4+gZMvuwd9lTy6Qr36TYgaxK8m/qQ29Y8lhtX5s7yu31dRVc3McWP7Jd6YcJIRjA56XFs+u
JfYLA32ZlFSVTbvE/zK6CiwiHbFQXZ74ajCNUrgpiSbpG80D550wrj+GB8a2b2JSExsOkftxp9k4
iAurqaa7FeZgaQh5NlDzzVHKAjtxkID+tIq7F5lE/XN0bLt9nG/SqBE75cG7FlUNntgiUP1xlfY8
xMtLnw26LLZweUwWNMrwAGwxgob6DXZtsIDIpEw6Ysg85z9L4PU99DqXE5PqI584SK1G4mqFTZHu
XBAd5geACQQdHqvoSh+6pDeai/sh/fanzKlWb/ZjTRZeUrZjF2Yn9/EJK2Khawa4wQIbur2jrb/A
c7MSyEiPnr5LZ9I52dKIaksgRgNx3A5d5pXhvd2qVm7zTa2Al7SrUFM/e7koT5xG9zVohDwEaOQL
CtC0CqHplD1BFOndBr/CXPvTHY4BdN6qsQOaIw3OuBseXnmFl1A4o99VXEWC1I60iuAs56bNWqQ2
2HKrf+xmJi9R51D6UVKdfyNTc3ux33B7W5Vma4xS8YNDTMBZPvxXhMwvvumlqOBypAGsdl/ZOjFs
0TCrEdtXDi1rUQ0oncv12InXtzqzh3LP1TntfIIZPXIjO2nU5id79yDRF5JDt7Cs9xoggKIQeX1y
/V4NFAnPywMT+w2CxGC4fK5ujhakdIF0YWA692+7fXs5ZoKGBYFNqtVGrSNPQsAr8zeku1dtR6IT
ptTTsCfziTF+MAK6xpexVRAy3FPPVQseU5S5BjoxYdxgQOnVK58+v92XGvITSQ1hkKQbZ1iZ1pSj
DXZRQ2fMbR1wATRj131DPrQjtqZUPfXj/V5GTIWSp9Jq7dzxqjXPQg4aeC78X81kDsypjVHfFOK9
/TDQXXyDBdFXrJmt09SKdTlvHTP3useF+AxiJkBGiC9aZqYh3ZaIrtTUpG5oQlo5DBc+pGxz1CWh
iF6G5vxkPqREOTg3euL4x0SjsxUV+M9IBE8nnlu9KzxhnQLScjkc046iBTvYU+4h3HLE1AlKOpIa
8DPBvxcOe++XLuTLh87+jAmv5oaMoWpdkhjC81wL5ZSkN2AWW0hEJLaoiJnMOvvzbY6QEaHYakxO
06H1CdgZHCPH5CcVY1WTT4kvsyQSqZzomqlSZSp3zxVAB9+Df+xDdZ6UqBEMlXE1z5B9UnBLED3g
3lV/r/7OrpLwJ1WnhiHQaJEZ5WCd20V0+aNLZMWJh4LOhUMMQktSocAOPq4hTYrty1jse0qN+zfo
KYmk/gzWdYPcnuwqq3Wwr3yWwhhDcT360LivrcyCAknENQdUziWA3mXSQEGnrl7pTk7MOt8u1qB/
epyEDyyVkpCoy/yn59ytyp/LMukTJGRjVBPZATkhmHCvGNfH28esoej78/3adL57UgzPZKRuPM19
mr5qf/OX4VUdbkmxo5HVtXiY1vnN123CkPxnvddQVnOxfjBTGtXRAu0C0PwDFEJeavtiFBHEI9dX
VoPqA62q/Py9TeaY2vUMelz9uezlQuv4wTabZOLp1MkP2bwCq9zHfOVdCNksjdU0Z4O3WoBA2Exk
so5r68wGux81PH2jeEcKQPN03MMJ8y0bVC7q+bWavnDXTr9R5hw+kesrWkwC6LDarmc3gxaSDHYe
JfUoP+mTaN4C0KZcUOIPMLoJT6z0R6WP6HKvEs1mqrO/7c6au0tn2PME+rLY1+nKJ1IEyA+MP5fl
UluVPHTAZDa/DBmEBL0I7GyH9PHRElvPaE65kTOoaq4fwMR/C7P/gaUy3TkfUnelldxYI7lalQn6
Umz+0cum0z4SL0Bg2JcMay8VRu0lMqxs1J1aoaoc+wV4SV+nnyWCyDZURSKQ06u1+YCwuKETsMwK
23wFEDeuR+8jB64PfhFfqhICoAZzmnK/RohKFjMyK9pq2VgZGUcKAvjeoaO4JVTd+yyHnyqyQjdB
s6npffrXyURgR3bVCQYncR5cU49M9S2CDkRWisXs0mV4noiyjMcm+9ysYdexiU59xgT1yNp/Xwtp
jr7eI//R7X09vkhSNk0lncGjg1SL7svi8TfkG6ywgywwA/2jj+pGbdlkSDIXW9PlFLz/2L2qZnGe
Z4XVKv8qW7I852EhHBrnfux6gTGSAcZGNjb8KluxfEkgR2JwEguSctB1dV5AmlouvKySf/+vGf0k
o3Ksy40QTddi6Gbcd0Thz/p8dEMXb6lLbLQTI6bMCNGDlKjFlbinGRKksU/iVb623FNxOC3NsDwD
058PlPz9JBIRJsVY3FNs/vtlyfIdm0dOisUvvq3axRDtXUiB0FTEGqxt0EtPqfBodk7/yvs4XJc1
GS/dEnNKsr17+kXAN/jWzdC3QOLwW2DL+wvlOKqyFwgF4uhP2skBaee5rGrqy3nwxmb/IOz/SWdz
ZxgzqAayfWxWr1zKdXDKR+0LGY04hCYXDdXSEdVpKMFSEpvCiDu90KX1sKC9Kk+UuDjwqBq3x7Rn
B37SyUThfKgB15TQLeQCJfCa2YIn76DSIu2fmOUJQoEG9/nMjCtp3WAirrX6ZnnWHZcMtPg0NpYI
HxDhE4nUsYqRs3Ks2FqIs/rpnoRcFX4VchthZR6smKFTLXJVJCQ5ZxWmDP2XZ6fgO9h9vfeuh7TV
XzXlq1I2dNDwu3jwjmwTgz1ukBHCIvqCckwyndDdwBxkWHI5Tx8eutOa9Kia4b7k0p8rR3FhM9Bj
YtfHsbTD0JuB5taySlRf+COLScr6W12NUmnynoaNKttAcKxXURXDFamxQT2L08JYaXDiIyU4jSMZ
ragHEi0jNoSB/axq3owheMIszfbFbIKppQF+R2pwL2HhVaEp/zzLPXqtk2X5p4JgdcaezXZkOr1v
X84E+H7ZxWvM5WDpddO1LZafYpW3CovCQrgENYyeCClr919VRa+zbnYbpbqdUGX5l5tsDhZp5WpZ
KORDGlBw3Exkb8GOdxnxB8FinjrVkggdo4vNOdDa/IFaCtn9nfIfY+4Qp9Bamt+MRFrGBm2+N2wn
1QVwxFfx8jHkMPg6SrUUqSeDnKq1VHHj2poBekDF79vEN8Pa4VdS1675q3GZntNxs0BmIcLe1af4
84YQQCGIlRAJRXUOZ15KNgRV0fsrMQg76MshKJu99JllDrXVKfiWt/cl+88ErDOGFYClrEFAHZO+
//Lhk6dSgnBnfgrN28y4ZGCnJEdeTUogqiEy3SIBKMQxoMRocbKineWMhrRHiwS/zSiUale/45GU
i6K36QZN4bo9O5DfEBPU7xU2zwsFUmPSqB/7Y9KMAyd9fiDOhWuomdhtbRzgELdK9RiFVW42Hxh7
YA3tQ+no8q5buHv3on8VAty+auDK3mataVq4rhYTSEzNhL9ydhefYrikixbuGzBWOvErq7c8IKqQ
we1S4FrORARavTkb55SSDqDWDiDh3EPzNkhwFjvKzFKCg1Enad7kbgDoKZVu/7MjeP2X5hI1BQmn
tGZE/2a08IVLMIa5CjhGtE0BWlpyiElC5gLMs3hBVlEsSldE+yY9bwGVhJiIiqAAvJbHui123sVZ
UgT1mEmT6XlLPgqOpCuBfgRoQbV5LPWQBHS74JD4QqtU8N/m1EzXru/35HJKdXMEEVWijpOR3rGy
O1n+obGFqY7ZArJzbyQ6FL7zwW3kdzK6bqyr3S8PEPSJTehg6OjvKYxiwhP5qzExM2acPHXLb7eR
uyatvO7Eg1APP0ygaz4BcX9VoX/kqfU8IBCK4Yf5wM8WDUMAvezvbYkgEdvPsA348nC/e1XKZDMo
sQAydOjBSMwThUoK8ygrX7QPYaRasv9eTz6FTfNzc10EUyj8ifFBRDT900rVsEdnUHb5YwS3vjYy
DajLBP/CVmhP2X1BR0T2FPBJKwsscmHoRWpWp9ppo6DBEn5L9MnjMDBp7gJWID9Rgnnw6GJY+5f8
EERgGsniip4yrbWAfxaXsB6BosdSuVW2kSUqE/khrv5mXkYRfh5qKMVYgNc74122Ny0EphNGGRIO
KKoMCXiseOlTADXIgPZjoThnqAAtiKUeMsVC1Xuq5ekkSJBhI188jYQ6kV6yhfSBB47cLJ/WXg2G
KSIwSmtHvUrFh5O5rdtlwxArEP3AdEJBo4MvcrqWlhO0+uTe40HfnGDNkgFupRq1qiC1ngNyEI0p
9Axm8NvWNPgkPJx7MEKAArsEdDtlfDkDdCnlcg49b9boFC2EsxMENIxpuau/pu4hkrcl9/lMowZL
7wImKlutaUZxuuqshi1WgvYpPILJBnUdS00c+Wh0LlaPShbXYb0VVSOAiiPsmegTKN5fN0cEec/d
TCcglA1d2cG+Rct9Gn3KJP+mq89/aRlMJOoVc9c6kEplGr7/cgsZ2Ujb5uSylT8kXrGP5PaAZLYr
mkDO5dpQnI6lESLY2A7h7y0+DHFp0c14JA/RFEf5DQ6uXk/A9D+QjF/yfGz3mBI2L3jjJRp/E6pL
VylvGF9E9F6U2Vvdpmz70Hcxg/DAUC5w/iJEwJiwyFQf2lObwEzIVr2OKuTxSj2dFEagNm624+Tt
c0Yo4fiuL9YLg7bDPZW6GwU7LdsUGzKdA6aheGUvAyvUuRwsUq2TUXqvJ6RQ5Zz5oSI27BOhoy0E
RqHx3thKwwR++qLAPzO62kf42jCf+WuroSobIv0MNro9mISZWcMB95bIGcMGRCnXg2BXzLHUes1T
mdSyvQcw7JT2PZwC1IExFKg0qA91UEwDgLzmHVRU/+2HCRqi5YJbTbBwM/B+MWAYlHURH8e5FbTL
xmnJYmvvHUbkij4u0s3msROT2RAO/PXI81qPCatOX6RS04fBnKqLRpa2lWnBbLTOmJu1EWqX7bYr
024HhJYvW6nl5SLiEe8ZtB+J481fU17ajOjT91oOes6ph3boPNv+oXa8ksUJIHfqIttMONCrOeoV
16xDXSualopsVh0Jr+ay7Rgv0EeLqfHf2Khjg+IZhxKFrBWg3MeCYAFQlGZV6uZ4UX5PnVPTCP4w
4p4MXQMXiQEh2De5bTGAXunlzToIiy7764jQMcmul9l6vfwXK2ed5ZYxvjlf3bVA1g3TVek6HkPR
Ab0ZyPVRtBeeLhgJgRxT523Dt/RxQr8EXTeltAc6fTwvSQfLasoSyWmueFh5+RpVdb9scEIiT7MR
bHNgD+mzMMoMvuWpmjac4/ABuzB63n762qJDIo/INlTZCKrEI7aQvrf18QjrJvpjieyp6g6uOSLR
JTmjffSV2LPdnTfEGnj+sJDaPiwKTzNwQgUrrVKr4z1uUcUPN93pfXXgtZTQkUIm2bepGVj0o//n
uvuPdsr2lmLtos9Y9ZkI5mlPxPSLe1ya694inu9uDNGKZWZbBbAYTCKB3NQL35tpdluzqvJfrV+c
5JjmIh0hlsDFssF6zjOzyzKo7PXwl6bShHqPH51p1mwLpHVkOkQCN8NsQbverxl1TXcy/WveAV5z
E0k0ZQ46CVbxpopaOTD3b4eo1QNQ18H1cwLPInytXtVSwOmfBBHggYAgGMf3mj42YDmHY8/ZZy8g
2031v8Kt7FCWTN/kpGJyO08WiMfcC+O8Bt/9GDeGAwFSWkAYvbkoxryaURY5J/prj/MWBLVVSssc
GVzrFXBWh6OHXCQBwLvxiF7V+Z7wzmxz6zLjGR5qfrgFWe5OS7sLmPs9eTuDpx3R1ETn6IoOQdC0
KIwYsxeUTZlfHWL7tJo/ZbYlr2KhSuajwJlTmI/ySYXz57WaNcUQgIr8Tfn4R8+Relug64JmNgwg
TmVJX1UsVWLNznQ7TWbD4i78oWn6iktamee+pVdJRXP0nS1HQLtJYiIeHVMqt5w1mWptXanJ1Nur
tljPWI2Isz4HTf1sB1rabNTAg+qtfi5GagJrHyqgs+xyPJHPrZimosZhiGp+UrrEp5cqy0i9EKX6
py53k0iPJoZYTL+mc/2jDLYEy125PMeU0Z6D+qnZXoj5RuPb+9SQC3bRH292p02m70IbvKxCUbja
MkrseYNkDTvNvBCRzbrPr1YEsVDzeyB3uWpPz9/ZuVNU6fovKGRN4I4SVV44frfTyhO7CmbBzN74
3LQg0/mWL7e5WnXRL2HqQWOPhPiOX5YgFbg27Y/EJiCunHqTqwSKrHxYeXZolrxZBOjnEbcqpO88
KcYJLcd2qe8laq8z1IpND6LeTfYEJ8r9H2DxmrWalPWbODyqDAWMiJwrks4PiNrPbL1A2u+vI4zU
yOgy5hK1HyLU108GpAx0fL7o1K5digVjIQv4gsFG7ZdYR3Vpb/RdbWXwwzP7Dj9nvqs/fhxlqsl3
ZwYEgzupIIe9saIjfgy5ZYYuEP0tx3GBBEVODyJVs63Mn81VV9H1dvn0pbg/G8K7MkE+gH6GPoyL
MoW11bOqQijLDlM00I8Zn5hB2WmxXkfSmhaio4R3gaA1ntgjr2cmyQPHyhEuaKsfeDQnrUohwURB
i+Hn84SAA2LVHXjnrSFUeDq831xf4ic7Fvx+VJXek8BSijgEqG0VGYnM6MKc4JNohKTKtIzrbnHw
5pWG1t4R3ttEsEAOPLkNlvHs9LBtOQXpD1xxVikvXwntNDw2CB9/OtvzK7TEHbLOuDIkxJoalkw2
P+ngLFNyCWGWUglO/mcRkiZhaIyKGR/mewkB9gEJDIGyR5DEAIw64nroKQZVTZ0evakpUgeN8P8E
HjmREtNXMGNWfgQY4xpdEd1jPm/FJUnirizEHAsYvKVc9Sqtwa49n1leSC5ktiIDBg3D13ITTxT7
Cfwo1OI1R/IMz325q/CXRj8UEHZrbRmU0Hx2pwzK6kivLjSgN85lwKhV5q4zUrFiqAumxFR0d0qS
tlmzLh/le8tsY0sPhOOT3UsaKPb0HVB6pt7V3YEfqoEjhuCnDRz8pQxT5xCF9z5811UQwveXCgdF
U9rBFunBP+MS1GwJmJg+zmap72IJMvwhcdN+Btf2grR4YaWjLX1twjp17o0LPtTKHpb0d+KnPI7N
Hsz8anf+1sJxkgb1XPwmlV8NqZqX21dOxTDPAL7cWe9ugPM9ADLkW48OfPv/FVn12cxj0UV0fzEq
wyJ5j0cHmrnzI+oVGgUVwA0WwsFauvnhcNpKBjX1N46RjPLmF64IV7t+jhZvAtcWJCyeIFnHTS7j
9ZWIXAK/7TCzbgOs5JTNz/zkgBVF2ixsoJLQQ5t8pwAEezZjxvnIjHYK4x8Hxs0lRLk6+3bfIu6X
Ds2QFgyYxEUcDa0crLYqgdmk7KsRgiQsnDXP4Pqw4jfeCCpE6gf2UWGbs+SPnCwxB2galzuGrajx
xX0z0g9ScR3OncEpraT1SlAmCzHdufvtfmXnYnIkskvJv52tLGM8+JvOWGyJ60OaFxYaIitmIAQC
c1q+FBeueyLkC6KmU1STL8QpQEDrDTCDP/rZH7LWr1g4evNGWarT2yFvJ3m7dNVix9wWUefss9U2
IJnVAaUjgHMY4a2Pj1mRMxGQKzvua0xErVKackMhdU7w8KpVppLxB4E1C4bFPeeQ8F7S0nHil34Z
JIn+vNQJoakxm5prgSTnDRMJhsNDqgO7hjIKq1J6R51tZv2R5YcK34j6mbJCuVili/LFLmvTHHL7
PqV2Tz+9k5sifUPEJh8ka4SYRsN5UVsW5fdKJ3dhCC1sNzqU61cIMj7hz03FHww9rAnhWlEyPlt8
5L7g77Op6x+QnmYAwBmwPz8PLQWJr3rR4JsQ0PUIxf1T8xR36ZhsmTkSIz6C6mIj4m0CLKu3gEiB
gI2huC98Tnn+srhql8IutvQX10m+NWIsQ+XtXuqJz1a2U6zm73YMcHnXAUEuH4Ulqx4rldehfRVq
gg9lhqLgMtrYMaqIHX7El8FIX7j+HHH+jYfA5I8FncUjo81XJU0aPnvXWV15ou4LvFtsM2DQ6yzS
qKbzbrDg8dajE0iRu0HaygwPyCzDCvgD66w2eppAKE0W7kMBC2195Ii/Ncb2zssO81N/uPGFFezD
dFcReObldghAGx5TiqmDI2NPOOuKAlDVNx+fchUTdZeXzftz9Mp4FCh7MmZdd1WizMPkGkpKhXOG
xUxgmVHEHPFfzCOFDsk4k31BXHT+igtIVwHEgOz2MAR7ATZKZ28f8qYuXK0tyle6riShs8CTO4A2
3CHQMkjmwVbjv7pUXnKUjhmhT8xcxzxNo/v1ImniOeb3DBPiEOMoZDCFyYgqhg/Fh8ulJiSCZcYH
DyGLCs0d1plvSG90GeLyBX9PGth11jyPw19qsr0aAFABDSlKcYaUUcoYSh7JCnSlHJ2hKPX886a2
tsbCsoIm3PdaJQwqriuJApr0X4DNqAXN6BvDw4eg7Ag5CEUDh/xpvP2W5siJM5IiqHByAByovTqM
MHuqQZjl2vz3qi/g5GRrzCL/DBr1cIttigxZxpDHCyIZ6+z94Mli/Dup+csdwwAY1Xc0uN2FR53D
sI89hdMG4ITnZFZ+aawwwjFA0CSiiAsUbq4/nRGW8vq7iYH0SgEEP3E2TmeTAUvlPdJgVS+qpLo5
Re7yw9VqV7uHTWyXPdFPyod0KgoWVC7I+mQg89q+17kIVUWeecUkEsUHwWKJCJqw61OYfQDIvMQ9
tc1vdGzclN+MkR3/O5Nr2Gdt0X+xELOncE0RRgF9wceiLzdc/IlqE3n8CrYjRSjnRUa5jOhZyr/u
khKf/FqP3Quyh/s3W4knWi7V1hAoIF9WivrCwJ2ANVcJYcrNGUtM2I905J68tf7m4MXqt+MBS8GW
qlI6C0rt/IWUE12OCD4Eh1ldeqk5WJ+Joa85LLExN/o/t096o7IXIBvmhajXPPtA8Vipg6/hJM3E
4VJIwIK2XfOSZJOu9t1KWN6UJ8Hva5CJegfWzSD2FTKvCHXIEBu4vymMXA51NFgXpinjMpld7PSX
cT7uoui9+TK7mNBL51at97SKHzRWpolNsxEbkhRShfXXkgpO1+r1gpmdKWKSh/b2WyB1hpB02bRY
TSHK8srKF16Pi4RlSHPhf1a4rgaAl0GRCfkNN+VobozcGgLVVIck0DKi/Rv4UDPlCbhmIIhDvBh3
bpZSzhWJo9VvSwtHf9nMWciIm1KUWvLQZlb7f3ETc1CYl52cnrmx93ZW0NQeNHuaNDOHY2r4lATl
Fiv6oA/kip/9czVVW68Brbc+s8bRHdQRMTK6TxCMUBa3a/ijVtRZxfFBZ+fQVo5hYxqq/BQJj+DM
EpPKUBVGRml46zSH3IElBEAe0ZosB3XXUwe0X5wsaShpKR6EMtAmTZfI/DR2rWdAq5uDlvBqgMBL
dFlVpQ1FGfQLurV4VC199/ZZud0JzHEW4K49tr/syV0X1uIaQkaQY8d5DWECs809bh8IKgkyPzaZ
kACDSbzBmH6kxALirR35I1mHZV/zfwx5UKz0jZV4NdOBBaHu4sYzEZo6N6AQk6CTtzEKTYtu8FDR
ITQncREXe5LS0fIcC+VJqQG14xj7OBsCwjN2PYwYSKGpTrmedr+EVevWroUWXRXI/jTu8j2QKdNC
SpsdnW1t8l9loawatTzY8JO3Iy/YKFnXITpUvcTPFiCi/8J20/MoK7QwCyEOJ9N2vcjV7D5j3Dd/
NTYrfES67gfxiTEQCOWnfZbMrm466y2bP9PoI0DA2Jse/3GG+yJ/xbtzNGXdF+y++Xd48h33qZnX
bQ/XqRSxlen6CFmXcv62E2BiM+7nxwbKs1hUtdRcw9/zpK6zr3xm6di8BuO14gYVUJLfVWhWFDrP
EZFas07TbsZ0apnHMWJ9FZJRZh1MwKh8UYfAy82eNY+hTh+Z08Ftw6CtLLgQLUystSwITASDQ0Ba
jhVxvVG85uC7JadVUOIv5CzQBnrcesi6PaaF6s13Tibysr7A+9hnoFsXhTgGj7QOeDFJ6C6UxgaJ
0FX1uoCqCshjrErdh5zBl81pfdc5fWlAcQCMkgQf5Eqcf+5ejq6midZQA4KGSuslruDyyCVbLcKT
egTTZZMEmelUk/mn/K6mUki4Zu/PsvzeCnxKkHFHKx9+UfA54ckztLJzG8Rnq9acQKSPWCRJ0WG9
nowSaJazccX/qmTroaA46dT+M03a9gywwUwY+N8go09LYOMSmk/1c7i2yIXlmh2aSNhH2RJ5nXZb
NFodbxGUwELk2hwNNNzPpFx1iSE1pr5FBVnyW+vaz4fZ9e3GdJQ3u/ISa5fjse+C7kQ/BAjvChom
HBBDsBW/MzCYjRqk7R8rAwDsKVuXgZu8KwGBSWDpydks78uy4ztAiiVM3Z5aEaUK9ziIHK1E4diI
SsHk2vPLMge043JjE4d1AcmjBbzMdqtFsfx853LWnmhWu5plVvfSAZq9bUudPp3zxPcgFmZQLmNF
3yFxBKa7vchk0M5urm0FT+4UsU5LDFOyu4dH1MSMnrNNR7NRxY28F2mvtKAcqTAdDO0tL1lOL9ln
YdZLZl6Y0sJGp8+u4VrWpyClHycEvzCOvA5cGFyglUArl2AKhFS9xl3MpszQQ730Ol/AY68Oxmm1
F3B4IWzAst4l8/SJgjaGZLtapulr2RIQwHGpnYyJDH7gjtykn5cKal8cZyizdm4HozXHMj02A6m/
5qIHcNIzH3eqo2NIG5K5lKjTq+R4ziNpCDlpvkUkVlNkE6m5nAX3OzhbgcFqMfxyaXfBTgJdEiBR
SogujulFthrpMWsXtxwiaxqinJIEmZUPYlTVMQKrhVPZo3O8WK4ZDIsJcD2cl3PMzM/fHTlnUh0J
xQlmvFGiD1tPVNexQ4rM60EgjART3QCqZwJqouRS53iPqmE+REg1hnASqB6gKGGOYILktL6kmuL+
n/Qd5DXzzwuALhp5tfksCEkFsK5KauaiBc0NKMyLPerWlQLCMd1kwHY6h8qgOlDymg1xY4WWcQyV
+Emonnkp7lYhvmTwK51HJ9333B3U9f2xnQHQwOFhyJhAeu7ucpzppQsuUFaiygdBhdegi4T6pCkV
/n7xHwq+D/nPK0GbdCxKiILGQn+PmNg96/36rGfBbC2e8HnVUYsFWEOs154c/N7PSDuKCQTXDCVi
O/uqdONiNGgdLshDQ2S3wwiC9/IIIIyQxKLinXiohQczb0vfC9uHBZ9SVhnWQAXnU7rTbtqNtfbj
gIt48gG8as24SOs0bgyjyU/HS4ylHWl/p4sWjQaBylV3FYbM6F70HLSgy4hlVsi53o32O2w9dfBi
aIJgyrlfij9cup/y46KFGJMC36OPkvuOKJ0jgkqZ4jqFRd7/lLa4E5PgsEApX/Bm3gu6enUi+Z0x
89hV/uHVdgs3dtlk7eiVVkilPZohILe5plDZz0eELvBnUkjHygkSs70wLignI/xhbQCquf7Jc6Pf
KIQ+pXveP2he6s/FTopDypwhaM6+d9e+SWpPQwKcq5PxWbiuLSwPJVdz6M4YiqJbl6Qf3NyAuOD7
aoyZlTKtW9ngPZ24k+nSwyuMgnQJUvEnzbAdpzHd+w7xJGe0tIGCNk8y2WQ+2/OYSNACXHJ2m/Vd
rnzWCcjLMAmcvs2Pyzhy0n55LnIIq03GoHDqvAp2FcRjcGWttYaFE40CnhRWO6dYik1pXuJW4M75
D+SoHgz0SBk8tCILrJa4yx/6TP8b5ISFmUXb1FE+a187d4n12swKwadHnUjTmSP/AlIDq2jE01YN
1wrVgtqX35BToZq80XqaORl9FM0wNxyseU5Bed8T/GfV6AeNmYC5R6xNznIuIR2dQ8iiMNLHSrMG
a1jozVtlJIdJc/Iv7XXSmR5DBqEgD8CATYl/D8iB2Dq+DFdg3PPjjs7rnll0Ecu+JiiKftpbrW4n
jpScFdNFVxI0kb+sVo4omGcZzvMgdJduJ2CYnbIyjcELPxRtWgC9rNzX5uuaJxzV4eUfp+DSc/lR
SALQxUxjE6gb+4YBQHe51SYVqLIaSwkyR3Gn3O6AAnwz/mMw1Lt7uufK/1UsybJoyMYpKL7334NW
aFcfUaX23iEnhcXuQrFd9ImyfbA7Laa+n0YFRSZRRj7IWEIfix64mJBu/oQtUfoinQ1x0ByNaaU0
+KwHVfot7huqui0H5QQMRv5xZvQMCJl9NULXYcIhdCU1nSry635GTBpRnL8zw4IV8n+q0w4E01eD
BnoRkOuxPPBJUXb8DHN2keSpsyGnMkQXo2U9kTYB05EWCk0Q6y5wG0TOUQGgjRkZtjL48bIDHCG9
VRxR55dXDTetCeQudH7oDyHIR3UxbLj8lcDA+eQpkx988w5CFEbhcdpUy90ZNnlBlKOL94uXFcal
LHlymre0BtIBQyjvIk/VxrD+qvoZZyJAHyVOUJtXbAVD8J5Qn7ubwkdoAyqBhXiQ0xdpoeof61e5
FTw5qWDGBeVUQfdmF19zPyqe/UVOIBzJEB8GnkpCceX8SbnQ63rF94TZU6rBuzcRblJv46eERX8H
zXpIS0w2tBxc39+KnEHkYVUj+clcIeBPREQOIIJJ3c9xzog0TExQdMarFsAzgu9qilgVo0YlY/cc
c+d6nv2Dr/AfdiFjp3Ysx3G84ZYA4WvjXSYQKlXY72Cwgnmn4u98BF1/TxEQ9Lj0lg6uN6m+VAcP
1YhnAW9yZhIz8rQmr7uiB4mBXrFriOND7hiy8bx4BUHM/4mNV30qHPf6O30zmb9Wohfz/08K1x4e
mMqT+LI2DFulAg+FLikicPd79AeL4Oyid83f8cO26LjqOQe+ZRjci0bALJDSxOoznJKuPvor2oNN
7amF0E1BOtO1XmGwV1rgyGaB8QcVq+kAZRwsGHZyw27c/PTUgIEHAJImAjDLgebNIgIuzy0x69G4
jX4LO9exIY00NnEG/SKhRAP4FdczQBh2b1Q85mfGJqrszVWcphPbM9U2sXGYBO+lqfWbzEPYbfcj
RK+nCdjDSyo/p/U8Qq/NKOmGfPflNjbGP6Y7FEDWzsfMPCsTxNcMS7oS74+N1WARnNZ1lD/dB0E7
ZH0kCvDieFgzAhTsH1fEqsLxWpn8x8uR7NNXNgmnetG3yo1dSmJ/03jviknMLjPfHhI6UtBGJgTD
MsB3un1AAMnfNb2oCcIzyEuv0QK/Yfovc5yaeVja4dJTgRDDs4o+/Cyqb6aWeor1z49H3UFkp+fN
JPVJYmnFW045Wj0QkgfovNdLpmXvahUV0k+3RN1H73fnrU+/hYTKqPFD9p7Ho5EnO2EvpZvSWR4R
caUYdQ6qz5oBhnwDLr1dTWdtN0L2aEBgDKk+cRdYUHuiPD6UNbBcTuzt3YaTaoBgTFe0lb01mT88
wOQjWImNkxAkK8heFfV1goi0nkZ8HeRn7qPYtEUrHB8Ec/W2DJ3nG4i4bUASC7NQHMXHegU1X2Ja
VEOl1grYZ4ZoDXNSEYbI9CnEXooVNYsCi+KRSkNHbcm9xle/Bn9ro0KPP2jsdcFGbyBhjJYYIgAX
a9TDVVq5FLng72368G4ZEde1el6mg99C7V3q5Y9Kw+7Cj7TS/XD5SfbJk4GQPxWIlPdMJ/nL3iFA
CJOi4baaUvG7E5k9uYrBFRraoYjpvy2/4+9Yn3Zxzy+OEvqq6TOn11FGm2D8QLVt4xW9qWlaBasQ
iOHrm1zQf2naAlYXjQfwX3avuzzhwkY4WS/FuaxtH65legcZYUbWb+JoqoM6Y3LjxGrfjzsJ3DE5
b/Q54CXJVV4rb+PhgHbL1H6WRIZXTNJMm2kcjRXqfR3+a/xxxJFtPF5vh58k6tfoSmvSiL0S4W2Q
jaBUvuqEqhpCrYrNpYggRSbSfpxAhWBNtBRNqWtBGvCl2Oq9undnk/zDN6ttWEOJS/WpWPuPEDFY
hd8FrPTw28fq/dkBD1aCfcdW5paysuo4RNRiRVPR1Gtz0bre9Avz5p0oREPDTz7xrM8foyAiDIz5
8501odXE2h1cUgebQrs5RmLQkolTDS7GGiYfMEv95++WLoOcy40/v/3s0VOuEQH24pg12DCiXYo9
mPteBtMVNNcQyQy6AmMJolg0d16+Cx+2qJIN7OUgesDZxz4z9CXGWq3l8xB8QszdEqjGw/VCxyZE
p9yQmcPaRTtpVxGH/64wFhoB14neiA/E8CL14wyXUtFJUHoYIAqZxS1/vAVa3IbvKZAEB9LqN2f+
PoBJPzb2NnXvuf2eUDTNYoqCj+VlreUJM69QCvrMkYvz8xD9dxHYxX1OWjsTLkqsKKeM1fhkj1rH
N750Bn5oeqq852f+TRBe2tuLLFC11mhCyWL0RxdT8oWM8KLP+wDYyl788siwZvtagMJb4hOiN8jP
76DtNtmpOrYQcxKSCpsj5Fw2HVAedyk8cJBQ6IiooT09wrBJMN9wHXvK89nqb587ya83/B08/nRd
ajD3qtTh4H9Y6/dhbqFUh1msNTK3sj/f7qdAsZPLxrJPWe2b6uaGbDtDObOJ7exlBBLuWhNW8lGz
X1iz6/tt71DvBgtiU2PCr9QSPDSF6yXhlf33TGFE8PfGk+AJg6ydxFhz/i9GF36vnt7cu6jaDA1x
tI4ujuRGqjwV22QCleyZ5MQIfbZb6wznjoO8kQOkabi/AZF+1aQm8It3m7VeHVy9PoNEIXOtnujO
J4Ua8UWhqcS6/cTI9N6NacDdQWNNaL9O3FM3z3YBGxF4XvQEF0Xt/2nhyfygpR/iX8ogw/g5Yn4Y
aFiJWBbvmT5l1b9+Yu03J7Zmlz2Kh6eiyb4yj6WQ96fONqbSewQiQ91PtiVasFqfQzIql6ZZY0YV
SWkpSI7YQLrEJlkhw5ARpY3Uw2uWPn3fwOdIYBiytZW+E3MTFnVJBYMIaL8widgWJVjBHpgeM3dc
lgYqoOfwU/c79ERU2uoUwr2w3EPw8LIH+V5H+zgmXMr/1JRR5SRyYoqZbvcjsF81noXESClqJRLE
mj828UI57epWa5ZH9b06s6CMGD1Zd7QGhkUJyNdI8ojI6uF5stJc4H3lJM8qn0xU0+Rl5J23FTnG
Jn8GEgB9q0Ty8xSucAQGpkvNindFKWvGbGD7ME3+6mjLRtwwM1RpmdJKOOxYSEkulpjeTiX6NKbB
WBOZS3MhOOnbYZp7f+vn/hk+KxT8USfALyZI+zFhf8WTizpkkh89flMydjrFO9MzO7DvXw0JENMc
IcrIif8PFawlBgMOi+VWk8oLm+CAkPBu+NCpWDaD++bFUhV+i5dTV8ZP+Jr+YkRl4n3b0q/derAc
6qNpmO38kMdOLupLAkre4kIFvK3Wah2i/Hhu6qRz1axTCZ7odJRbV4NivQAJ2ulx24SXNpvBfE/L
5wCNEmD1m2oubM09iNcVZxma/RRQTOKpYl88ej2NKWc3B8qeT7oVMw0eRfat8pLaX4qmTMUT16P4
DcmPxODN7BJSF5wmD8RaRFwgEKMm4C5o46Re2wyhkvId/49iN3WfT1cx6ojtEjZVoZHDB6m80oYP
PbDx02vo0vms+ve/VNhmrddY4yPV2pjzqILLKwlaOS5rwK6/PIl5M+Rg1ztIJOzwiGsjt6oLgRpq
uTNGErBwLnAas5ktKzXS5PHELnqmTqpKBMGuUQs4KWUh23YYXeQEa+1ojfMwnyi+05xj31o5vQc+
uhfB9weGMdD6zaF/hh5+Gm/LnytAFHZMHGgpuoC0b1O5Nps8Fcu93wo1qX7Dph/dvPm4X48djOxr
lpNF0oLylIx31+L5I8vpjBzcw0bC+iy/1UWrTpNOlBV1Ry7rdgEHIemAmmT/vCn+ETwY6lgzDL18
E1QhSRfsmCsOaW/CBNVa/DwWIX6735/OctkeB7R4CttAl1oBvdPooXEXeLsxDtrn3K48qwhs3RY8
udzAPojCU5WF1GrnZp3+SJ6stHtQWDp5OWLitBkL9XCOdXLwhPXReh9HyobpD/f4D6YXdwRM6Gq4
N2U6HxslGZwxpjXDUh1qrWW78cw77poVymFTymbKELoM3i2MAIy/3uohSz+UwoGRrjBJAjtHr3KK
S0aDJJ23MyZK1ijsu/KInI4vJWT2sV2TnW2rY8myyokUIbWO1ysBYLaZf25YnpbC1zAGOTafNhlX
Qw/wZou1vVb+5S1YUWuLRId3UoEDCVATQWEplWK3mUqSQxmF+avgSRRjkODriUThFBRgIo9fyiai
nRHsWpssc2h4lXnxTX+120vbkb3F81HeK5GllpnFvJuY1ms64ImXukkUz3XmIdbg/dT31cl4qHll
727zc+JMDhKpGZtMy13we5GN6DRvTdjqdOSvtASRoyi+9R+xtOTRFVAATaJw1ilZraw3guqifhkU
SISrW/6n1pQfyfsABjtKBXdnmy5gVcpJqbzUpW72wyj7ejC+ltZGJ9p5+nkayoHTBM9aw0v0lbbF
IY0w5RdLC9tHVCCNRXR1nE6K6xfgqRu2eMYuNmWC2SP2VmglnU6IIgnl0MmgqcirZ7zB5i/QPI/G
EIQLn0M8EDb4sjH5Umk1aNIjOjCzlvD0ssT6mUc6PrqSPp2TfiuQDen5yq1jwar7J81np/lqokM+
8vVJCa60/mnehPLrcGj2Bew3pY0aRaX9KvAudskKgfH5WisMbku6iqEE7UP4zRxeFPcqfOROhXph
s+GAYNiOF7coELw59M5xbYWCYZeHVsaFgLAYgBL+40vB+fcQfCJ2/L2VQNmgnzCyXNv8W/gz6tKF
4akhmeUHGV3Qlzz0TVRPJvkfo5/jXFBXuNjKav1ZZQZL8hb3eLTw33QW+pgMXOArYXcl2z9eiqGg
sf6OfxFY/jA4s5FSqDV86eEi+JVxR3oh85nusSEFAh7gSiTK6DZu7e05sinbtCYXe810B0BEoxdW
AipK7dxtBvIrToWifyJrCa02jtvH9gkJIB330xSb5oZ3l/WHrtozt+wSt30Eh0bGPnKkmqxZ/bcv
YjhZHUwx4D6mwRnk62yPW4YrcXungTK2FKgz38UimURF5GTtrW6Mqu5a2jyt3JhxdlOBvdfvpSLd
wzr1FZe5Q2EnmvbWurRh4a9NU4KAitcRQD7ecmh4r3Ui9itZqvC32vfaN5kNMUPV/QI++OxOYSE4
alTgZbrsxrHZ54ld7oDaf/322PDtaKEd+JNSyaaqwjvsZ253J3qzETk+iKPbxE8cJYdjaLtta0Vl
/hXxgDEwwTfiwLM4BLBZVklellJOYGtSm4/fP5INqwSitY/BFkACNTNFAumZ2oPAbeJyf58zfw+j
Yq86HHPA0JSOu3Cb+/7xX+riGDjwEb2v/KiyUwm/4d130zmarH1fN8vlyWanlHX13Q+ZSsBuImfk
gsZTw8SFpZZCNfGT8j5r/HZVB/6q1lR24l5KUeRzc86FgJw/W8WJ/eCtXUJ0UQ8NKIRquROQyoJV
iGovm1xH7tLKEnrHUx/FP1+9/3K1/TpiX0NnJbXTT9yq6czeaLK3scfNpYmSQk0iGKNNfaPBppE9
m7HNSl2JR4L8KK3z6sMXoHsldiDGQ++rBHW/zzy/fAwEgrkKsNLTZtjT38GPpNdFcGJRCiRPEISr
qr1sQfuPuZ3/RtlA9Y9mNJLPvbhx5sK9ZDr4dYpLVvMXiPs5IOWIaOILvcXE8EHLlks4VduoCkBN
tDthEABxrnfw6pJQgM25u69iirxLZfoolwgR+wXA6zCt46FAhZTR1XXg8LtM1lhXP1kfSF5YzbjD
DS018yvorP8wHkNmG/v3KEiCL7LzQE5C/yQnLQ3Ae7aj/0x8jVwyWAQlMrPa8wzmTt7ww2RK0bk8
y4qjR4WgoQFkhVDjXbfK47ylKWpCpYBogpMPyceeItOc5HMmzajJ5UZzafqUHQCHY5Qfr+1QrEGj
BymxUrhESsQCbv73UbcVIYi6NcpLmo8wrCiVkUdFKb3D8Tdi3BWB8bC6dxW2r/XAtkBfDtH+8Fmc
RwQS+EW3HmSQjaE1yc3J4HNiq9mEMIKplsyZN1ZZMoUnL+7oKTUf+ZLQ+k3WnsLW5ZS6zmx6S8ry
aoyDzm0j1nB6/8zPKWkY8DM6UndKxX0hGwNNLYYKc68/nkrMa3xHauMoBQbjSq3OSU9UqWqpxRL6
fsSaAtaXvcM9N6dVEbsYWX0aWv0nUwWViuCEpgLV0SILKoW+fug9WBBRCfSK4CQrLzrqgDXntCHF
jGVFKPJYIuyQXuZulf0IbWhuAyIHrDLxVLQv4Tqlt/Mb0V74YFDfxRjcXFU71PPl/+SaabVgmibh
Fk1hYd8rUDBfltBa+GqKyJ5q2QKjvmRMtd5diG+R92H0nsYRXBEqidVLe6JnmdbZbvr5sEnakCIw
CnhieZArahID7yqjSeiM0yhanI9ScuGUKKxqFWpetpTQ7DqSfvvakbasQjYlgcOQfS3bHt3uSEyE
Zr193x1+JFImNkxcT/DugoZqEaRyrmOBT0uZ74jzk2404L5Af8JfOn3Hla20gJTYyP0DP2HsQKM6
hHPEKno9AX21zAJTAo7LhZVB/iXLpEs3uBhbIbQLP83cQceSImT8QS7aNGp3sx0SnDqBE6XdUGdI
vGU0BL3pfDtX6RoClfUAKPHDnGGTYM98lknutNpu+Uxk6x96YqGVUf77hNyqzJA4nDXAWg0Nmj49
vImA/JbH+parGVwYkNRqxUI0EZcUnsaweTQ2tnd9O1HdY8M5fMx7dyZAaGSP3f/uPKOtxTa4R2f1
R/C2c7gOWqzfDz5kC5/UNxDT6zZQEf+5kJED/9bFv7WLoMhg/L4+PqfJqIcGxcczqDlLZci+9FY+
1JcX2Er2Vyxysq1FJ+sNjWLJ4gZu2dhY8tV3rWqFmRYTOlsq7FQ+tcDqpiisb8sd5EjlpPGPcGD8
oYzIGZQbpa6ahHlGvKWc4WcsCBEP6LQ7ApSGw1iP1RS1lXeSXt0l5R1ZVH4QqX2zf3684VnMuDfh
yZj7MRCFsP+p2aCqntQyHVYKiVFLFgFvY5w8OyiONzMtCmjiDX4Xc9oUhCrLLxtYKo9qaZBZAzXd
1M6zdSTBt1eVcCXtoBjGxHyrhUJGEK4+RgbAdNtjeF3ga5uTu+MmR/TnqZZrZ0R+t8y4cavF0cuj
f5QYMGYlCHFk4gfQpjGQtK3TWMmnTzzCF/RMA2HO31hOJYztOJ/hFBuCG9txkIX4Ywga4fp+2pqB
Ic7AXyA+ywjTPz2WUwsVgoSkZCl2RHowS2Mdd4ibav5u/2/EWkLpvgnounUE9v92reL8NOJaPKt9
N684eqdm7cAUXsyZX9Z27gEdHZwQJgayotHzgfzVwq6dBrF7bQ3EvjJ9lP86e1UtTTL7RZdLuqHS
vEp1usXuzKMqPInnKS0rZPM+iPiuew1xhNDzvV0B9Wvhu5FisMuz/tWtRtqxbSwfy78fXogLII9z
hclS44uxa/2ED7VaIcHUt9rhynh22dL3tztoxF7uMRta9r9VL8Fca+s3zqihfwAWtG6xoEZJ8l/G
MlO+gxilM3H8KiyE/0GwIfgo6VQHrz0SSdZ7MX/3tiv/te+ky4d3mnaftALbGjO3caK+ykxEsdmm
jxhVjUtyhq0TybBF/jbfNBoKpKHFsKjmLIWBesJFlJr7y5pf1uQii1nij0HBS3P6yTBJITRaAb0r
28UZnll2GDLPt1l/DOJJwp35Zel0bf6gNC+d/bb/EsR68gi5SQJDyuaEIRTv9xBKQ5JsuRDnG+YA
C/UF50xteQXEOErnSSzGIjpUCOJroUwN22DcaN29JY56AXYQoJaEYm+SgzSfWjaBZoURGFjtyN0+
cyoV/UAICV9tk6b6pN7Dg7fvAxhHIIi58XeJ6Eh7mFq7qK+Uq3kED+eNldxIiIaegBlAyPJ4SwzF
iFkVGb/i4Gw8TMITa7BCN6oLrHJE/eebf08g1MVDC44tMj48A6vmB6l3BYgeICGN7umlruhQxHkH
Q8wsPbe1zD2d5ZLCJxduESmIUAtbWHmjXnH/GYPjZcv5XDrXYtW898cnn+tuw+pDbqVeF9jjczsr
tsXAMvQ6Oq33nfqARVJgX9GeThAp+3onAmXm7UtjqWIMBkyAmN6o1Jbzqtom0/DVwd36acWmQIhR
3KhwH+uYtYE6urFTFn7pHOyeQTALd9OlPlGVjCXQds1PcJDbwb9rNwNiEkLtXLmqy2xm3H4/Veq7
HDE4Gc/nBfCcBQzHE5sktR0BV0JfKv5lxcinyGsXZQcXwRzaMn8GDnkHO+DsjSHI+y/+QazPvanI
72pcL+68hTCJ5ft0iGsNJawXFBlAld7p2+XrJPVZXV9vqEsOOtRPO3Kfkdkv8PG8ND0x4CKaOT8j
iGVM7mAD1U53PwZnXuaG3IMQsCC/8HU7tPwVFgwZwprdbdHykq6MQ6V5xWLcgohTrzPdwpiTrph/
tfQBETTv6U6yamiIM7HP4VUQJVnIHv81oA5mjyoVTj/juIYU8nDOelyLC0y+2pyVXimgGR6dhBlT
axwPhNI5m63LTYljyAEFupxwMTN6zWdDDzw1oXeicJUvXYxyaMmdr2NxZ1NZX0e9u53RXGcfmjtP
5y1V8JKqB9xtKt/Bp5FTJ/AAHqaHtKoTFlAos981l7P8DYHMaD96sNBnxOvOBmbrlrVFKraTcoNN
o7OsW1Jzv/Uv3Q1rQYlmlrYKS6pfnMZ0g3xSmQohAyG5H5FlmxIDuvmGmBJbWARAUSPNRjd3fMbT
3XPv/kMk4vWRE0YBi1hWGYqihEmNmMNyeNaAegRwFn4FKR7IqH2ONZFPBVgtQxYmALctgE0C2EYN
5NMklvnud5+6w+fdBjDKTpBaF7q6iqTsXqJjZ6IoCmyvcB9jbfUEr1V3LlrmNRX0WjSQJMRLZwgg
DZ5XLHq7vLG6ujYAp69EwOkG+pp2rv+HWiq3wAgtH1KZtvZ1E0HAr7s4pgs0pYrUhlN6VSj+cUKW
dHqH7ikSj/GD+X3pI16pIkmqAwpOoIY8gFF7Z1obfxE/XndlqLFh1tTnSMf+RsaO/uehZI82jKMS
AgfeRcrrrpY4YikprG7y3BQzhMEt2ogeQkR+wVrWUQDCSG/nWPV0kIkbbFcZIwAc/ZEgjVBcal/k
e+HQ+ULaX2kV+D1Q0BrZIPFYQ/YeFW4MdlMF1tuy2Ip2zzMK/qrhXBqRjcXjN4qXBQN9uQcF8MI6
96vSYPgd1SPejVhfxy+8SJxPbKujPuHio23t8q9carqYighiC2mJs2u8T2eps5bnax6MWmRA6Ykg
rE4ShvX5U58LRhv758jPHn4uipqLcpuFswB3zM5wLo10bHVvTZbge6CvwvbpeipoNc8u+G10vmzU
mjo8X7zcvfpVpC9gqxGrb2Ycu//cc6V62q3U+MEaR/AxNFYb/Xl81ZSJdLkkk/7MjLbvSs0aV84e
f3VTwn24ORNaBVU5dqM6MGgPdcIDkZLTSbmWYS2X5GRbHnRCmsziYvvZSDR2l3T5VsD/Mi2hfm8y
oTgNMVNTNlWLaPqreb8AVsqW9ENauw4zzjucJpFGNv3uiqURhio41NsZ2qvQgY5arKU52bbIqlya
lqFAvBpbFPUvXe7Z/vWHyWIRlRe5uKbMo8k94eDhFhMi2BocdcPuYIj7on2ZHMzsQhDKHos+CHpn
MtLejPpKInrindxSAYKdifBzZJH7bghN6CRYdUPjxjO/t7UBaztxe97J669/IhIIS9zBxdsOEAB9
eEDEpQiB2h4sOPCPZ6C1ltAv3MHVY+AoAHLmA9aDiGPmk3PIjuEiuFNMbA2EZTbMEfn4KpKptHZt
iBnW7YUs4I9cEWaBC7ISFwUUbJ6hCQn/NI6kH3wSX2YuoPUqO+Rrj2twm54sZvRz/q4vgnbwBQJJ
6uL2ThpwYK6BU4cewDpOE90dNgvLrv7luNP/2WLkNc+MMYlTJ7UlTqycMnSwdxVBnts0Hp8xaQdf
rzfOcgAmiEZMBabigponEmerVm303WsTxh8etM+RkdpBiWFw5cxVXcKUEEXddsbl0Y5MvB/d0OFl
DP5h4yIEbN2MDgEmdLy/hrdeqJZOqsQLbL/in5ZYMh3pXoQGZIj852ZnejVybeykegInX+9c/o9o
/DV6/Z+dtspD605roplzfqCLTjTFO8HGd0+ivxHfnzq/k3uGOVCGw/6GnJP6Lq9668a5Z6XZjtjC
4tCaFtsibKEOsMJfIYMNHAxn1mTyDvE9FpF27jMmmw8griF6EXqgXqXGD1urtfBavXLp6Xc0p+U0
RGgdl5SXsTtFZyKyS9KQhtr4O+3drsNa9RGLMi2Z/2/94Q3tHmhD5OcOGeYFjQqtjQLiHO/znY2p
BOe8kbPHrCL3u26B8ATr33vnHj/3Y49mASbxrDqygLCJltMMCNuxDRivDy1LFKDaF/hAHuOdIzD8
3ql0W9BJLctS4h7TpspZ+RPFo3zWHEco0slZb8NZZeA4s1jagBiUj6w7i/Dr3A3hsf5gtmK6Y5ck
kCFaiZhLP3mKyo2udjnLNIisvnLPti0vGHVTZhLdDJWUXzb9t3S0KMfkRaJbfghPToMwBF77czm9
429PVA/RzIUWgtJP0gEVVpzur23ecNdY4OhqTECOzQaTlDW+Jhv8AXdHgrpAeozPwXTTB0F1qXgj
hY8bisj9WdNYKZtZrqblfnxXvB1q4OOA9a4+4ID+p/BGHvx9uA2745kjuYjPL41rhzJNb6XVWt3g
c4oK0aR6TG5sWdgkEn0Otb1+jBbM6BLdLRhcKwi/kZELL/7o9IFmjCmADCRgGPcgqqOmVPHXP/bJ
GJKk6G496UtT86JqWfYuyqEEP5q+G+fiSswFiq/iC8aqNn5QFpkkRcq4Alq/8IKubGAws6x6byOC
jWrTlz+XcNg6z7K0a7jWL9HFoLwxCBbwRsSg1mqMIc/RtWJCm60sFbcz65DTX9/GdldxI07yBDAm
Zpkpgj0ExZjr9qzzB6Lkwhq/HIiv9eUC+IEOTPGSIvq8HmoLchgJX2ZMlgqfEkpkGtAB24Cb9ExP
3UxlkEyH5bV58KtHZAbMSlPPGZqUKENZ9VWSwfbNya8Ti8vnFraPC8LHQ3b9bhpitcEiasvFjS7B
UIGSYRTNzajEQONjXP2XWqhjaMNrOaQv97NV4XJBe7BkTZ9Ep8r3i0sxspOvBrnhknc2lii8OOhR
0Jlsdds8HPhdi2bFQLjm7sWLCPcQCjBEDsWIkOgIpYP5pHhs5aIoEY5yXQIRCIuOF1Z0UE4R2JND
FvphYdk8hFHawAlbGc2qoAyYilXvShzhnTPsd9Q7Ig1xMGh4fYmtNnUljRXteTFIJQBHhNgsMh/9
e37fNU4bIMMVD1fyPtVp/HvRT2ESF4ZahDntvR/ytCtDByc1jypl/BfKY03PNJagTQzKnoagXD05
lBNAtbK5sJkk3YEQnMwqjdadQHJpAl/K7mK4F1y99UWMybZ1g2zwpdFmxaYx997Sq+JWQYjrr1mz
FoHME1o4AK5OM1PzzzkQMAlpGrTtCjNbReSVwuG7paP2gevcIePEMZvqJO+BdwSHRcbjaVwN053S
chsoc46CZNXwZIb9SgL4RexXP8lP03vBDZ8u9CZq/vOCFQ6HUEWIRroRMvqE72hOqAAFtoinWnw4
Er119SgQ/D3K25BUOrVxzGBOAUi9p/a65QTHHpsXZRSwqBZP1NmwewPg4jmQHhiBuheF9r5bJsUi
p4Kc2injhqELxM4of5pA4AX+CFllTiogQYsknEVjvYSI3bBb33qerKRbhGh1NNbWd6Pl8XTz5Ntj
pm6O0aRRxPAL8tHgIKTtCckeSqDcFCjKdT5iD+BZqJs9xX3O681AQXm4VZ4twwv0CvPlPwjd15Mx
hl6yvoYEQ8SZ6NRo0/RtyXcpnTw3YbVlZEXapmdhbUTSs9Jqtu3+zaEJig+d5XRpiAsjZMwttGzb
DEPNA/zY+CfC1b2Dl6TDLHPcTd6HxLLv3ZqA7hNhy2EQbSyH7O+9rj/ltGTvTZxPq/NW4H9WGEKn
gU8PYM4CIMAB6Pp7IERMmcWq09MLzCEBVNV1u4cufxI+fvew7VdmxypZaWOcC0u27hVSLtNQemQi
O/6TiL8VQoPCMv9RhCH0l7CoNmFEcnPdkIy6hvNK8GbCeZTAmOlAAJehPrgBLk0jelmXpglDT4rg
KtwB1asQjIriQFPSViHPJTeKmOXazO2Cx5HNp7XfibedQa27y6Y2tXsVMUlmqKJ/4ajmqbO86cEx
S3yY3pXWCVJ+ll4oE1cyS4RTDsCyHNAK64g4Ajwbkl6bGFZZDqZLEn+KP65IqejR1fsNDj2+8577
Jd4gDJ/bCHgvHyifxeZ5YTNsXSwGHuBorAMvyEjc+NNjxhBDmsI4dLeA0RPuZebzbfod2Lmwpxto
6k6WURCfe3sV6UtWEjVlM5qPMU+6obJbxXbZpwMrZWtVDITWoBPoqA/GSpJqPgt9r+h1HBo9rHmR
Dqi7arNyCilL+uVE7h1renHxYdQks7oQ68nJ3MkA42p7mjsXWdKerMwwgJsDKXH5fJYx5w67IFVD
c5SPF5dwzQonRdtV9oH4GhCAAdG0hGnNIxxzW3s+K6rIztANqkWUlqQCmid4mhqiBD58dn7TQPP3
KyfKzzEBM83OaAql2/0+IsOI0eL15aumxVybjDrpOgGxhjCGtEApRKSXx/lVGv+5mQGfiD60ZO1r
R1laDZV+rMquEMwAZMx2ZFC0R6X31Ca8B4sN9PBoW64wL0AepiJQZzNcGJ6FyhNI4TZrOIYrXHLl
1S1Fll8g5pij1uq343b0CRkb325gBBHSXWInxilyp6yQMRm6KWRdgnp8UFk8X2psEg+FqGO4GpLa
ulSdrwnYAbuw7rckzCo8wxrtsNCzjNvr7RX9l/uQ9Gv7SrzcMR6xz5DVnZ4D1DjY6CSlfTpn4/gL
Z8/f9uTtt4ntS8wQe33yPpI01ZnYtD/4cnrqu7wB19+XwmlJHpOMNyTJa0kziGCXXtZJ5gp9JJrc
zBk5yDELaIoJp+MKk2Hk7fTmKb0tdeMpD6BFTWgRN2a+9nArjXC7wzPp1nkPOjOXP5+dM+QkqTq9
vBxh3dGsvTy0iFkwBQaf2lmsW9VAqR5RhF89wH3Qub9myP4JPgPPwFiSwiXCCWYiKT2sIDRIUKAU
F6STQL6IWdr2W6PiA18JZjPF3cvmfSiXgx+vWZojXyYInqNK5FkcyhKP1XmS91UihacKTjnP3ERH
I9hkwPKjv1V7N0j0531p+J9hsgijdvkAiCSL7IhqrB0JHqfHFAPjuHA1tKmlhjd0C4iEoFSLnTbL
rf8TDVeGHjR3E35KjH9JYnRAOudvrlMj/m+hNO2RLIOxiupFPC8Irkc/J9YghfH84dlweid3suIA
vNq3/0UqrEo0Jpb7PjJj+w33DDUVMBic1yo/zCElOeBn6N92+2PhIHJG+00QOffjg9Sn7pbtMUci
RzAMo4Kc0DxoYlOvpenGzaIBEwH0OK7E3sfpKJIWXUqx2PlNIr8e/tzWWDcBgPyM23leXOgV9Utf
jDhBRSjZE+rTdRlXezbk1Q/xxygdtEYSffUlpWC+9Uj/QFsP0w/xWi65ZYsEYuxtoppwWCcTUfVv
1YZLFdmeFR/NmpJAsDynTKMbO8TkM6JbSN1ZWH57fhTU3CZkJG6oTLrBpsLjW7Hj6jTZ+ujdSRKc
zR3vYon6EvW7VAZon5v2ju2vmVw4eFYGS5c1+fc22D85nsHqyxyFfXc9KodZQLfEXZ8b4GXEVIUs
vafpZBF05R4RVOE1ySLShX2xkkuSPp67LqbGAV1MKjk4UnTQ7wiCqE5FjWr/j+dw+0ahbW6WRn+8
EHQCJhPZL1aToNqEGNlZCfSMAu94OEGuAno5MAobtwLKZ/Y/kNRzy1kuZIB6rBJzGkFDD2LFGWCa
ZcKhNTL+yfx8MyYZa0spgKb9o5ARnEk+R5sDBNKQLg5EjqOpTP9H7jhrmR7ZbdfR7T536/ht8zDA
n9DW8LcdVNGagmbpsBray/s4oy2ZN4tDqr2BIGudJ4MtYNLI5W1tgfg4IJRYecBadMjxnnIU21/7
e8EbSUUBh/2QIvhnI60dG+2+IFktQDAZt6/Z+AcmDGYXz/fK8vMeIAzNx/W5JIU79BYYGAUeoPYH
Rv7exD+96eQdDOfT1Cc56v1jNa4bqoxJZEHAjP/aYc/YqS3JFRx0CJo+3HACMayDCyBbrrfWp0uV
pfemxdgiY+Eqx9y3WwYWH+8zayO7UN+iAIMygHQH5OeKrdEoM5wav0gcvjHAXY5VFwXO0eGKFbcf
3OZF2WXSNXRxQYVAuL1AV2b68q5MtgqHHrEW/4so1uvKDmijQayrZLQ7nMU1Mk3I6Jj/p7MblSyE
etLEO6+ndM2YaG6zTRqiZhl5X6n/dgSVq3/FyjGKZzHjCg2CKkdr3Gym1GO2B7A4K9tkR4YMT+kA
q36SdXqIzW92YyX9KfdgsF1JoTE8QD8aEyLUW/KHIZpEjWoDeYSb6IoTtt4mfCuSfmUxQkqs2YHQ
pbjV0lOVIr7H5vsN3WBc0t9OWKGUkgoE7ZjvOEqmrzuMqVMktBXgzjEuhGSq/nfILQsWhYIbcP4N
7MR8qykXl8jaUEDDEAWM6kZzFJp7JAI1I/Fe2q66opf9lGfngIXT+Dd668pr5k4nSBPATQNZzYMA
oA9gvq6lisESOOjkuYvgmt+VhpRtHskDqHl9PvliZn7DV703WxzQUO+v9x2mbncdJyjLYFsHRSN5
bDqbqzDVYW91vs8lQMBIiQQxOy9odxSIYdFCguFcUFrpmyGaf2p7SEtInUC43jpV/uv9McEk/6UG
TVvDlARrxdQYqcXr+AZFOZE608iAxhsVEysbmTMwqSk3F1ZU0Av0/r+qCAuTpwMH2BUbOxQJRplQ
h6W88qHo81f7sDzUK6KNXdrEBUPIVU6xYxGvaj+vdqopwniv6SRtnsm/sNVrhSDSPnM1uP+DYqS6
ejZHZqfrfudfK7w9G2uXtPiyUlpWcT0XjW3Sq5byJGi7l/fn5UznzXjidSdD21hZ+aqMcJnygW8q
Ol2bp3MJiF2rxVk9cxbzSmrAh5k7b11gRwbTycb9xxSZHx+yhlLQYdP9xooI9vccPQ2AyqEHR30U
6tovov+L8OYgP0JwUUhNZXyg1x7PyGxNgbUEqr0LrMRoWm9Al5uiMES4PSnp7AAPh/lJkH3aBng9
ei6ZKVM9FbKb7VE6khLkJojoldiyCwpduq5HehfG2bAR5D1JO7Y5catCzN4sAzuJYUqkszYBfIfM
9ZGF6R+vTAMwfyqe8ceOcS1opQgVMb7OLrhSiSWxdcw/qwG/So/p0/6HvebWPVIpuxCVrgC5shwR
wRmXLrrFtIAbYiZa+Z7XP6l5aChu7iu6nXJLi80F/vKkUnIby62SI2gmdt5TazF/gYa4K41j1PrO
+cvuHJ6q797a+XQ8yKO44vEpP2kb38aHhdQ7wNGWX0L18ObfCuPa46t3xyaHH7CtTKtLTVNKVTeF
vMCJUecBQ/XFu5Pw4OlIgmoYWDKr8HA0AEjPsD/N/V4c89kBn3jD7Y4i720rQiU04UhXI+ZLMHx3
MB7dMRk6lawRgVf7NRi421gc4GlJKVda0842aKMOx0IsPSt2WoBmn1s0Bs2id8aCGSdY58PaoqV1
HUk9zZOOqnHtfCWy+H15kfqLyyymR9C8XUv34YcrWHWLCAWejutAwErnk4S0/oSFYlZMCTVl9a/m
F53SkqkNVo8V/qpUilzuWJ1MiJ22ZZKicyKGtjPVLc2RDwqQWCfCU4o2zzMtB1ssvJHVPnIZrUp0
GgsgJl5keCRnEu+Omlaa8oE1+xePcFeDdCWDfTvGOf0/e4VJOzlY0IZjUUWLF9yMmobo9d7FcZjC
TeoXHAYKeg5dCOjnUaN1g7oedOcYe1It1Va3rlMtYUnUghDWhgDhIWYiR9dBnylQUR+ipxp4WeSj
XbghZ42woYRu4sxjqTnNxdqTliGCVtKplHwlgvMAgVJGkWd/+R1RGjWT80+ZzfJnulv/dGpmH08R
3s5dbi+0OLwFCTc6wJVerZ+fUeLQ52XSkXowTVwDjzWkjonBuhS9jHBF7omsfIP8T2Fc+EJxMhIo
c6D3jSW8E9pK3E7Mz+rh3yAt4QtLJtVkkViCBtCh3GagScDlhZrLgi9a43MVAbkxrxuZM+Ykf9/h
dFukCU2mgMJgmlAPswFcrDldfTcDe4+l6AjpoVpeMRsfCrnUaST9fsgY/kyOcHU+Y8G8NvebYPot
T9Su4JC3Un6lLsRSc+Vh5nXHw6WxHxTwOCnrpqjH4wmrxOGNEvyh9QEZx9RMEiiOfg+qp4QJBqRU
C4BD1wtkzzOWuOdAdcLHi8jL47w44sUrDr2kwthLqdIhxcijJV7ZChGfh4+QSjb7Q6hCJd2ScYLR
gmunU+VO3ZmTIeW178/jAIPv51FqPKSUU/MU1BSE5LLBRsKHpSEppn5eS7TWi0/cmp0VrC4gckzY
mVmup2sE5eGtbS05NP44bXvYxcMojijxkERxqMNNDbOnl8/7f+C+3hX7aYtAKvpIahfASUraVCom
/5/xrcY3zFS9VumCY8ma8SybOikdG3R05xjhsOjTlFkbbGIpKaVwmJuI22RHLn9Tq4I8qx1gIWdg
NHmoY3/WNJ6vqvewMHCKoUCHZ5KQKEplg55/8AS6y6U/cRAMUALbkTuaPtaEat/hHUyk0n6ytAwX
FfVj61s052VuTooflpH9gbe3GLCToiS60nBDOiE0ay35oirMR0voxMEpHRytJrS3YNUsdLphmWTP
FgqfpjnPPmkiifLa/hDj78WfRJ4b8GQQ1Lqkoy8p29gz6zCDNTUyd44CGhI733nCm9Frw1A1wslI
59spEyguiquS0c5JNW5q2jA/NT0A/FSdY6Ye9+ZSstm1oS5ml/vvFl6DFqiQcFkoq1a2LmLBJWd8
hSqEbnEi9SOxXbU99wQnwPnKSbqrSgU03zGy6frpzbiWAlaloARbEpQjsfKlGlxXxM02TdLF87Vr
hMtX6NCd/zUiZhyTSo+o2wNTn9IbXk5KLEbB8I2IK4MeW3CQRhKwmM+ILXMtbY3dlWrrwUIVF947
QIEkGjUnr0RqeijDave1kPdLkH7bGL7fkR9Gn8Px04s/AvWIJlXFYWZDqyDen8Dr/QQzi1V6Sgnk
hSmJFF5NxJKsS8wmcpKE6j6LISD0nzX9poOdmgOprER1jmLm/rLhSiraD12Jq8ZfccHDoKQUJ1q5
dO3uCH6eYdoG1Rs6yeLPqcxPxA8ZcSLbGKjRLQthx49e80uIzXWRcU0CQb7oa9KJu3TBfdZaySpV
VuFqOW5qmgCkN1ku173vkTi/jevfOI0lgUKtjBcfkPWRzZDXvbvLvh86GfIJg6RQr9lbQmxlxldz
R/ZBNYaLJTUJkzpDcOdNwy+NKsjs2wXygKeorCVA3IR7ZekJmftAu0htzKcqyiayCiN+AlfD0/hR
IZSSpDK51TbSrqNEUt5w6+ONalq1+oiZQxJEdIst1qvp12bjtrvHv6mD0StvYikPEX2W9F6LufkD
YVBs3fm2GrrkkHJxJmGLLkUdMdFe7OT8f+SrqL+biI6Sy/3e9Qo2HXZg7g5UNr3mUzETqULxjzjS
VBHjf49MqMFpVzJIyaAF7/TvW1mBqZIxuNVTTNkRewavu3gdPJXPdgbaxjzDsfhujoJBRBXiTy8M
Kcs8j+l9v1FMcJr8MCs488u716i0Ua1CHYqSKTm7dIlWn4/meFt/VeWwrYEFbRQkxm7Z7e50zT9D
oKRFZHJz4o6nLUKmXmHFeJPG9GtNGZbjwIQNozVuWljhBn3IHmUI1EIQrI8ZX3hKLLti89p0jAsD
xoSJ12rV0ffoug6aryciLEEclxK3S760cZqg0/yHstgwFUX0YDsZf9JvmSkAplq/NvC8x0UvpkEJ
leuYxOySbm9+OL/L4T2Y0/eOebMzCkc5PQj8B/r54184eTeDtPgwPeZhiDvC/1EMtSJMRiMBQj70
tU7Ye+rMcW2cYkEnQ0/Y1crfxUumQtavB53FFmyd3CazomscozQMpmBm1Te9527ETE94fm1DDGP2
bfduq3SroSHh/ZfxzytPQqZ2mtQDL+ZiyiB4zDQCWvAMFhrt0WgZOreEK12sqRwF4MmK3ps6CL/8
LbV1964wvho2XlfYPosI6oZG+B3HvTzc8vmZFEZbP34OwmHXPuso6cdePZShNkUTNV/pYewEUo5t
mG4V2sEhuRyQxpoKqtaBbihAzyheGEG8ga8AbmpMgqwMjlzi2a93KKMrCZxm18ckG2HPMMDCm+5d
Z0VQZP6FYtesijcJtX+Nm0Arbb2POZYEF2SryZlOns1kS50u1aqrLloeXUQCzU8/7KXCTde9jbTa
JOEeW7OPj1lNAUM+/qDK1px19GHOJ3tRRCOemXmxBOYcpSjS1HrkZl2+/KhQ1tM5Jzxifat4EupB
4RY4AZeael9al1JmXbmY8LG5IRILvan5NJf/5Oz+dpXY3ZVrmANGb4sNq/iGrtAnAY4d6Hyo2TQA
tU2ogUp+GJWAIUy6fi11CanoHNGRok+mIu5ijBphJ2InUO1EADbnRKAkwxHTCc1SGNrR+BPbz1IH
H8XVb7tGuNcLrLWaQ1tPpqIfjMW/5Y2aUqhXgboExTJ8ImXMf/0kM1q5Y/2YluLFcPrcpIeLNseX
xfbBAZbQ7D2j15hcl58aYGxPBe5Q9pf4c9f87IBy8HnJGR1A0xEYnfiMhltyO8mtnNAyvN7NEZIF
BPPY4yyeH8b1Nfr1Q0m0MD8vOBhEhAJcsNjI5Qne+ljepWQaxYlRDb/i7rhUV9+pk/tVk/BKWV5s
W7spJykwyld+piU6Wi8ZNtKgtYu3rnkiX7nhf4BfoYw3IlZ92pLSLhJLH3eJUlOzJZegVoschTH+
RFiKrFiOq/ykq90jM4UL4zJTP/Gwlt5D6EZcHtp5Uu1WFAVsIr0BjacgRvwLiEMsHcwGvswBXXWR
OMFdZTNmTegmRoik6qWJlyBKZdkH9j7ao99dC84mUc2IbM3ujimfWVV3zh96YYcwBBeWLF9hUQu8
kTrJLydCfEmgqwC/PjTGgq3+dlAyZROEXTvCDTloJVpJONL8AYNyt72Ue+ma/oCikD9+5O+dbxNs
7GxqN+QZGtcKYQiu6Vuqz4LMOXbIxAACwoaxGKX4k/+PaZm8S7QkK3IJnYydxlkg2rtJIy8p9ihs
bP1jDGlUFddNwnpI7dA8jZkCFfobmSFfD7n8kgzeltiIt0rXyX9pgA44RlyaSKnmK90OlTdJ6VQk
Eim6DyXVJfug/Wdcm2yF0m0Z08TLvtIyj0QHStYJUsx913jXFo/r/eZZaX8cE8uK4iHhfg6ah1QV
M57AP6oZkINW5JJ4fADXStIwAGr6vTi7Zw9qEPMcWaJrGt7dyRjnpgJZ8zP677rzTNP3W2ulegg9
t0vq8qX9ijQJnK1C5AqCf/SoZ2fhAvHR1ahP5lm1GyN4XrEci5kE9kzZTFg0biYo0LtAJkNaEF4O
8/UItXjaXivD4UK18B1Jo1GdoJ1e7bDOcuP8bnIYRzSjVWbisoOyBYiaUw+M5PcUML78ng9zg3pb
gP19ycNNWtbRG/YVPgpWVVV5uUFbU57+IOFyvwNhR/q/aEXhKMLIXC2L2VRNlorqaBPfuk+fk2Yz
p7lWHh7oNxpLXUMxQfewcc7v+2WnArSN0Sop0CFTSY9tP7VNw69ExNdlx+CSit/18CGqW4CPlEum
HH+q/7lPDAnTElY944usIvFmjexJYuxRFuN1y4sbRq2zBZ/nBtKTvRPzWJovMrCqVHiW60uc6Kkz
vGGWyPOsMI/QuBevg1ywlgunW37rtcoLIDQnQhRPCD6MNVNSgWo5FTYBhobJ0a87pf8KAMTxbmlX
x16/1vWqglNV+zagQStIO2eruoGfC1oYBj4lT/s/sy9uWJsm7DtTjnXokKhvrL+fkdN+BP+qvyS6
bE0+tCoAPz0rS7MVD1KJ/JSYMjIEdT72MOX+wuh+2C+VM6kVRpqb1LwgPE3H60MYxLUSyUsGDZsd
kyB+90K3qav+jieiIRHFj0bgs4pvq/VjJ7ekBYk8m7RO3MXGX7AuOyU30z/oIbLFSK6BBNbvQQJV
OlN9/sjSYsFJl1tlX7uwerwHuu8T6Vfwa6G17yFpKumlslPoTVtudqh2fgW6gY1tE0glp9xrav42
gP06O0LcWKjqft6/AGss5EQfoupbtG1E77tiwupFyGvIjFWQyBNI268FswAYR6VtfG80UpkCgqET
cDM6ySQmDMkpwG2ne/iuzIe49Pd0eyWRoBv+6FvnMHtboVhDPiGHxT6KA62jm1hJdfduForFSZ9F
dvIA482+GKapysh/U5gtWGNWsvcuUhvLJ+ZsVX0B1OU0y77VZ0ADwemT62X/C8+3g6c43S0CAESk
uiCA9bx4+3vrwDTifOr98eViISKNPgJuO3OOAbaUqxydAYmSlOOKs1pFxAaZGg7XIqS//C0lG4nv
EuqYqeFCejaZLVypdL7HGiyvegFyeM8Exg7Ro1Iwx8aphOw+NzVP94BH55ijabFKFwrmuyxObXi3
Xd0CUhqY55uzmQBFGnktuTIsDGgEnhmuOzeFuFh5yS3EePIiO49S2mW8GuaoWIeL3lIHzZGywtEX
yde2TxU4lB4XrN06MfSk5dOfVbQWzO7frhsAivWFMI8C8Gd5vzip6eXCrSue++GckthatmLBe4qp
fZTxfLEFGQOc1Qfjko6QA0885ZM1fDuunuMzBqgOr7CGFEDCmUnZ6o58JwJ9+epRgScj50nBNoZx
xjDZqD/6ZQYhJFBNof2OOaTbOHq0iHiM6fLYILfOQS3nF+LDZd+vjokAsThzoQ1bDbGi60WL1KXy
EW+CiA/mgK7+EP4lJL0GMRObzgMEcokwfMd0k9uqax7MlPvOippRmuY/hwEjSy4hOyI585cRv9bC
gkRFC4vzbo8POUhpX5jCIgW+a9WMC4pWoTXcFYSzwYves9Jj9JleGxXQDRHI4NEUIg2lM8V25fQe
2q2CVU6P4pur4ulhTYigr/uDnMwDex4oyuwdQgANlT+X1gRA1nMMksD14HVrbVyCQqJ4xbCSMFF5
fAt2+WznC6w/yPmkgW1BQ7aUY75U+5C7TWoOtqrianQEF9XwM1lpz2mHKAlmb20vqgR5WTQdZeyy
XVjiHHaFzxkRQ2m7t/bT4arVL+nA69DAqx03LFT/YuzA+wioXCIZn9zZ/IswAFdSjyKQsOVo5J6P
nzEj/MG0QIPi03kITg+gSre/0OBBbb5jUgVH7PdXM+e8/2IaJAW7DoiZ8zcvm5IGMWVlZBSpMpAN
X+0F5dMZsXk1XOvo5KfSKm7tMQCUKFLFh9RkP2uHCA/fU7ryY1rsIbeARONNd8uoArbnBym1c1Nt
QVJIZefvGWcxGK7NhItBebe9wKI9/yFp2I8QH2RfPLvtvwn0xmzqBkxa5LS1di/YnKnXv5aww7Or
fqiFbl3n5eTxOXeHcY1asX2R8UL5cIIxUSorYQwVq0WhvyoViFwvYfKSjzvWHK1MiZ2cdPbF05Xc
1H05YP16QBwYwExx0ard/y7MACCWpvX/BenCA3w9tVW9+CFc3s5EkqG5wQETv+nO2f+BGJ7zQpsL
guVhuz8yeZVn5CBlJTxt3XGklbDyBTd5j/Jry+ZlPjB4a+KGrZRPhfiuDOaDGIM9yjwk0cPuqvSo
jedP2mxUY7a8mInngb55/+Tau7YUlkW8B3eKbmYSWb39r4cNn4zM2z//36CMQLDrZcVJdk/lxEjU
1Q3saiXil8PslsCc773x7PGgPD3sy+98rXYcPqkGmNjKmhXWx0noTuE5VRqP6uiUZYw6kwdPf/NT
Brt8CjURJme3u1UWvwx2upbp/UMVJOWdjLwcD2IrJN9DjkbMhD2zjAce4oGQwgH88DuSNJfW5U1k
7+nRfqazw4K5lwrtvlOsOigGZV0jZaQIi+A8hl1kcJFe9a791MuKIPN12u4WLgrQKEzwercWYYHR
9LjzFobnZcVUgS+zwJg/jLCsADstFjWQFCfBoCSfBXCt+KQP6BgAwMY+0LF8rQSQtzucxZSeL8vq
2RH+3etLEfoAcCY/zlYl13ObtbcWYvwx1QPIbH7LE9ZBGOfG1AaZ9GRDjxeujNovbtlN1greSp/h
o6mpVybQh1ul55/4xSP3AS11E757LFXYbfijQ7j/dipljaom6mMTpwhIkmfF0U5ESb4m1PPWA4/Z
5tf3clCNYlHfdJXk1zb1eTbhXecTeBjtU5TmsYTjA9Ww59UbKNftS8jHcdf8CszbAZkWWkbcIrQO
0pvRPRFW5Xp9ODyLM1g4LhNuv/ZKkutbAHdxVs8CoxO0Hc4TLzuCYomGMAu0JYqxZoOHJWhYjkDB
yKI3CCvtAKk7y+gMIsF9y4w8fli5yiGrrVg434y6NjMzBg8goFE6G0zpjgEHn5wytG3MriYQZJZJ
Wp/yYke4LtoBPB1suCUzRimiGwviTLBoAodD0xKlrNqMhUmxbPxbjDFpsMc5pjT3QTEaW2Czpq7a
6kM/haMfVIP6uadc3JaCfbtjWvbETn0Ag8F35lbzint3n8QgshoYoV5f5MZGHKRNHyvA0DJL9i77
YeuEEZNxWGuzU0bVF6s2OEcZr4pwui4lBx1xXAWCe3EXaGVrNZQ4UcqfTdvVnzGoU8R5Zgx379FQ
zfnZd0EOZb2tNpLu06bAThJ/hdyxAVv2MpRE3mdIzJI4CvV/2sFUUXFeMeq1bfG598N9UUngO3Jp
7VrH7wFsir3QT6eYdjg/XCe6A/9NX7xcpP3IvoXlIoYTciRFu9tTXOvpno1Zmq+0m69BASk7x7dq
KWEKpyWQM2/2F5AMixhfAomgcMdG+shF/dfyPfgo9xGJNZ+oX7wm21N03ODzIduXUNwq6B6brPqB
m2+7mrjKJmLhuHEtFNUcspPsbNnMxPTq4SAA36vQ0u8/Ks6Cl1K4gQemy18yq2pBkVv1eL3P43+9
TRkQBSqOwk8ir/QXi0OGiHOFwyZds2LnOVNYZyxu6I99HyTSBU08edFtdo7AM/9hX+KsOSXxnAQx
/O7abjR6SHTE27Ike8TkDAunhTU9jeSgnt3H9PAgNDdlhzwJ8M9gju+IbqAO8N6HZXXlGaIimGW9
7mYk1ph36+JbXQaR/nrvr9ObtDAXLyoGpo3ma+XT4gLpPV+bekWpDsjuUAefRKq7mGY0idLoz7oz
7/Uf9gFI1l/e2vUr6jGFbaV1kGGnxBHVtMyyUV4V2tQhTHEj+OCPHrOzEFeX57oupoyUBsP/LrOy
ZyDxM2HZAm3qfBBCuB6ncTiMZHYW/hkra689IAdN96Dwe4GjVj0PNMteZM3AzCrnlldc9yoMLrMV
fUyiPMny+hJ0nWmz3GiiIloZoQlHxx0BT7GofarhfT+TxSWrW3CIfNev6PMS2eWuY3NdxR5dSbQM
MLIdLLGJwr54CT5VIAqMcxSBqzRptRWveYY0QFJq3mWQl/BptqbZNnWaVvYgVv9rnGSSbrwWo728
axl1x4+rKulU+2MNFvXRZGSlKd1l/IZuh5ugxeg9PFAfHZ/xD0HEcAxkI1yme2nNmcJIBI0vC8nK
Kj99ki3oAXnPA+7QRdDKOlLYYwglTMgpf5Ht7gVAauzy9j5udvGeFTRZs60IK94XD17wvRU2asMA
09wKjWE6gYfgwYbJ+Vt0mlPr3HmZ+PPcoKlfLGkLHrMMjSxJYjto0WTP2Ur3j1bqVhicblSYFRAb
WW4whX60AzU+sLUP2lJl1UeOAU9ObTpIS5R3hfUntJxusrlRomcTQ1TG9slhzq00HVwSCjlUBuc/
CJwTjTWxyhRR5Tse2xzfm210tQllXrKF5F0KAAlA/8eSja5d5H4qY8R/h3MF+TielPqF3PkbwpsT
ZLDOxFD3PP2bNq5QVEln1McOv+nUUViy0c4F55qhC8Y7IX/tE7spGXgv+Rc2zlz+XdWiI6DPdNDm
Pq8VN9Zj0q91qaibA/BeqoVdoZr7oltf2TlEz2ygHhSLebXUJOeMvKWIPd+XyZn+e3nFSyw0q9xp
mvinlMXdDw/01IYgwKejTVH8eGdAxHeuhQ1V2vY0szWFY3ekuQe//VTtMmT4ovSyAFejmDl74yUO
jS1LvlDBLxOb3I2A9484uMu4BkNkJ8wSz/wi2n/uX6ze/wq+vNoFqqXsjpyrfHpjIUtZZcjwNJt3
2V+0SxnHbyHZbTIcKyPXE+kpN5uR+Bn6CG/140S5/ZVJtv6lNJWY/56DvqR5mM0oAoS8cajcIgWU
w8ymLbW2MK2KJoC8bHpLW808cnt5YKrJjXGXDhveVdKKnpI1frZcuusf3J2cmsfyDv4W8Ymmln8Q
yzbP1zR0j1gPbYPq/i39VHxj2yvVB/vjo8uDdI7hDYGT1HuPzoolbSURnSyX3rMlvsi9+imM9qOx
v3zI6VueSiQR2doE4ml16zOIQ56qEEvoie+a/o6UdT8b+4ykD05twehJBJMDJ8/y8IX6yI90XvnQ
fpDk5J4u0Ndpoci/gPo5mBMLBN+TXPmRKmyu7FwYfYgaFbPkU0081lIUR90IWZeTywzonWo9/ull
Cdw2PuCw+q2cjTw0Ob7P0rb5AINz+Atoe/ROMiTfkDUU6Y+V47AEaKISLf50aFkWYpGSFu153XES
Hu5DU3hzjLlxcb55Eq9uj36NxtTn6GVR4a/H62USDd4nuVy4MTW7i22S3LKMYer2NGx8z5rEgFNW
RvkSBvg9zb6GPVR5O7d1zub4RZ2FPr88Hnmw593Glvd0kMQJa6UEJctG/ZCZ4RpQRyrzAJ1rKrb4
Imw9sTM3KP6uWWJD4pJdGEYNrnPAxN1jkwF/wAYWAG0vbAg38anFdAdtd8nBafk4Q3IK8Eiz8O8C
elaOaAItF1k5/munGCJJfB7ROssCJKafzyvp9uE2fa+OJfTorLqmeK6+jMRP3Y37/zi7E/sjAXvl
S1k1yFVO+hYWHru+oiYVrORQyqw966umW0ud05E8HK3VAJ57HiY1mbFJyKoJJ1E3ElHzuZn1n+k1
t3havkbjL1bYvubmztndLxVIvvUgzF/TytJtqcthqfu6+cHDhmJ11UWkhOPlYlVe8G+PWvEm9Zta
ENI6ld+nBoYnJy/SJ600DVZSO/Bkl+LJiEaJsoN0CzMTcv/WPzYyjSKWIdUckNXlQcY8UdSUVUOO
hBdYLu1ymGHXQJeNQVwBQynBU/DDmMN/P+TTNMmAEDrL98gNM5LGCijlLIS9UiPG0IGfEE4gTuh/
Wh7PxcRn2fGw0AFL1rpF9xom6nNP3MmrlTmXSNS68RMx9asF/FHMJUE7joJggOnMYLy5rMHPdcKp
X7Ju/icj/xR6IWPCdgXeBiIAXQHc1XUDoU38sSSFw6n0QExbu260l2SoJzChxZEr3stHDya10Wqu
LzoKXVRU7Atew6qV6CxfnZjujnYI+PeLvU93ZAh25lGzTGO1XZDrfQEcywrTFG9zl9XVYt1j3nbj
HNzXWkcKzj5Vnhe8dEnmKEMMozdZiH8dw+VCG7k5b5R6VD79J2trLevGk4lYut8Gmu8l9LBIKMEo
hRb861Hq4FeBBKMm7BNVkpK0uIP38GXfgMA6sq1qlwroNM5NGlnNHzHmjMw3hlegGU96G+nKS+Uo
Fx9bZ5Lgi4KBVJiFHtEXGPbZZ7/cc89kMl2jQb2U989EshTB1fs7zEy8DSWX+sF1TjDhPzrKw6+l
cArabxDqaUQAubA4k4Ofl33RrqxgHiBryPekl+5uZnBlrxBon/WzOlt+Y/NNLS0e5OVpV468igBc
+KX7GAABcz+9ahUxlpl/GjrtvrcD1h72ddxluFPBRhcDXIdG58k8tQSPPXNN0X/E/bpluKz4J7ka
NXP9rr803Vxk840zG+rbhl2Hfhr31eEVsUQG+9V7ZxezGQF/Ua5Bxt1H4azxlbMLR1OM5DMbVf7x
SoEwPKMvQ/lsrEjeGY8h/G1ZO6yV4eRk1eAk8yL0UscSmMmCYbaD49EvY0CV+sv1t/fNQHAItz2C
D3TInkQ8t1paYsCxzqKdkqMRxt9glEUrZKxB8lI4iXRrz5n8FvlkIXmAlYwkJOlRxXK45SySjGQ1
WHJrpxz0U19X+tEwYl6ESkhPiy/gmAzaRQMt0TC4W2HuinqnPuflGp16U6pHP615DdsQ6oGMuH1S
sIil5FTLSdPOl/zFVuqiVQdZzOxidnLRg0Qbw1SDHk4kxiW8qcYk7JW6wYDeZbKqJ05cAPX6OK7L
0FWk0fMjxgZoLjT9vbjSInagYyu9MxDjmP8IqRh+4+Hea8SR11CnZoQAwWZBgtU4k+IlXXLAHuWH
YUZI2xxJONaL+mYS3rYvsUfZnI7C0XmwI+UYKr4Z/zCUhafU1aRjk4dtREH9QhyoqFiKNkgpZ+du
E9IL1BK2j2bd6ytZQ5xBbYpdUkkdD59e5gzqKG8A/qJCZHq2ml5x6OXlMSK/zZTIdHlzEy6WpW4r
3PJ8lxbgHPrwlbRaA3QSntUacAre4ZWtU18ZUFtqo9HMahJsV63tZivn57g5GmjFhNeJQ7p5YMwF
NLk/EHCDro7oMMuPu7dgteB8bbdEtE2hL8Q4QF6JboLn05RiezgBeL2weFJK5F8RfHwi9mR5+QY2
Fi22ilWHJb12rR/3QckqMSY7ggOY+Dx5ogWroOqKjYCVQKYAJihPAGfYhrdjZBZbL7Q2/MU/xIU+
ocWn8uu2D9JVYQRvarEkpbx1oehqT/0dowoRAGTl/ikGziZLTpHfl1KRoqDgkCim/8DC6Fq/baZc
jCHDWh4UTvWyw2uLqk64UyphcjMKBvE6EBIQwGR4XfO/41Rs76c8MdfBIl37vmxknJj1O1uTcWGc
bbLu/X8X4wC9OXh+/HXnN7yyPOUOHpfSMXQv1mBBaXJVO5Vq3N8AMZDvnAoLPZZ7ItPc3BGh99ar
hS+O2qqRfKReX2yDDCBLgV5vMqclQ6h5lLoiiLAUmFNMt2xqkAGOAyHKdDmQJhc12MZDGPa6gCRU
BCe+raj4OeAOUUpocImsBPKllSOK2MrBi5SrC2Mg7PLV1namyH/yr4z0o4cZ9vqV20kC/iWRYlqH
MDOw5loSTbXVk8IV+PtoN6Md4/oOl30Qt2cJHEb1dhufm1d4T3VOdlcqbsL/ZNNP8NhNXiVEakWc
WgHh/kyc70vAIRKD3f2dDzUQ9vSQNyabilQZ2fcRtuCdm9MjmCPleaQeEBceszTUbTqfHCU+Oblp
dBKxSmKelgbrjSm1cW+U4N27yeUpxR4OTrKwv9i2yB5AL0MTkXtseHFeJDYTZB9gfKy63EsV2nSf
J6HyPqvCyjJhhfy77A9CGHppvELWLnhXiv09pjO/tDFl7zz6XzeSwcdKDPXHAM3nccrrG+9rE/Ef
dgpYynP0BElwRQLZF+iYUDOgYoJ3asi+8NRZ2nLEuCdrxgDzkk7fQ5GHUI6I4v+Jy94wag95xvso
8opAAILNf84DQhgKMTJM1aodZJv4jgcgnajsJ7mFNdql+qD2/3kOpTubsAIbzQRZyvZ7LhQMyt0v
k1+V5hk++Rk/7VEYtRbTBsVF/olEAFoLFmMoEnDUVnG2kkFaQNeo/xjK+mn8PUcmOTY8ZcwzT+O/
/oGeufN53XqTKxuF57L7Ben28FnIO3dO2XZa89p6f54TdV11zj/ghFdVdfwWGJGMQBHWcQHviiRc
ZZtpfp5jtdV9wETFTL3qXET+CkbVs7gjVIHWBJYV8Tcyyk0h5RgBaXi4spC4pNZVaCupFHaw90FR
vGYJmjNWzg7vOnxHpFR1vmzNJXUoPMt7yfRvcJyc6+Kyd43BHCOVVY/0/fklfSxQJP07MsWfrgW5
o2tmuHeSr6NhoKDaBD1uNKgY1l9DzfveUkBKEl6hi/kqibd6jqOkRt95Wn/ATw6l3RWw/gFHz7+o
lvLfEUNuPINy+KXGWYWHZ60LWLeUPVWp+JV80wv4u5u4C+9wykH/EGv4gGWHwni4MCMiPvqreFMP
jth5qi8JYSkYK9lAg4lm6C16TWSl5qjK+vRO5pv+NRB5qvYkf5rJwcYOkwip37pJaSzEf0cGkamk
UM8SvXRLkWXMx7bLq63GY1ytdY9uCpSJ9+hZ92yA233Njb/NNtUZo4yXufgSUvbFme5uc/i5WOFz
c2tP/F9tIFU9GtwZs4UJJzz1MfctDDU24O1IpwbO/RSp88NLdJX5Lltpel9s0hOuZWT00vEhUC1k
xZb/V7C7rDdkjKsDc5+APf6iolCpRYwmuOHbsa1C5cXLJp7+gMPcsYUgLxhQvLU2gWRhEU6AztUP
uQ9ryIZIxhwOiXiialSxg51ngTGQMwDA9iG92a9INx5xWkibik43Zn/hkda3BFvM+r1TN1dTT2Um
ywdd27PqpL6AAGxqjXQlppu5uTbKaPvazj3VA/KCqoVozk3qZfEg6dc0D1Apy4/fziefR+6IAMyU
2Nze9Ab7BuIrQ8iib8Dztpk2Ermn+t1p6pUVVhzg8V+BakyS4d8gAhPvSBKVMhrhTbO4mlTHRmBU
R5qm5jAQPq2mUJSeIIXaWDEu7mGn4BqtzZaOsUpv7HAJ9bcNmx13c7YscbvvspbePOTMfSQJ/to9
sLHRD1qJmPwBiPUirJA8bT/Bpx7k5H6C38IRpScy7GZUClkGjZs7t15iZVYxK2jp4eKppIlPAnPI
mT2UXxlFDhUYJAcful0zbkG7JjyiIXLMlpkTlOnrPQNm6tMnS0opVobFJYGXulE/+bKi7cygXaVc
OiheeyCHFByc/4vjjOlL0ezB8p3WJr/59gxWTcNgsPUWgW2uJbfX6pQ4O5BK0yFL+1+NM40JXUO/
aJBUVaFAtxZlqhfvZtKkv0z0e97WsSoZHfcwuIPl2iIUAHfJsXe77s4nKJtSjhTprw/Z8WR3dY0r
2i7VK7oZaj+jQlheXPXoFHB83SZS48vh62XCMSlHo5GSLaiPCyrUR3yRxo+RVhMYDWm0d4ovUTqz
caoicbIFQctsbWV5t8vM8JI3Cm0pSpUa91WWoAVKePCrGFHWhKizW2s40mkVS3NJ1ff3GaKQFf4s
R/PUeDAiIdBlAkZ/Wq0Fl6AHM3NjbhL5skMgYx+nLHUo8C6M9kaJ9CCa5aIACYWqHqSIIzZ9s7vJ
R9OfCi22+RlMQvrGxOK/vRUAKsCgRJ9vSPNYSJdDy12HedX7a0MCI9M+R9ZJg512UbdqdC60xljJ
s4o2BNu6/D/2qvEnGVzU84c0SRjQ5ZY0ydnewfLazkQ7zA63tbss41Wn6Qz4YTF5lwOwiMFJWE2i
a104W0tAfJoerZPxY8+7Pioopl9etZ8Hu40qac1arOqOsRESdhFr6q5gK4aIa1mFeNU6v5bytkzB
s/qaP2duSe9ZcSZyxeAWA+N20fKOfgqU0d7p3EbvwGLhn30/7AUsdQJMI/wvjW5fEL5dMYc7yRuS
e51iJTP6p8jDdE9JX8xC6DtRzpTRH6xwesqBKfWRDlYcnsfq7B8Wi9FVrOup4oQBd0nURdd8DFp0
F6wBCA1hTTLdYUcJLv1q4AY+FXpohi17aZK/iurwQwlSU3c02n8KX7l+pu5IDePVl9hVhLBxrrpR
km7bVkTvPWUNKlIjVwnu4/9lcoo1rnNEJrmvRhFfTzrJbIjNxjxL/UaiB4+e1vZVpoe//S9DhR9P
fs2yhbpYCrb7Ms5wQCw3AGO6sVz6ckMfUxNyfwNHy+7X072QNwDKTw2ZRupB7iDVx4Q27gWKwL1+
g/9fWfTGwegMnoBVU4Xo844vEZUwXsZ3WBzxTJpKvwS8QOyL7hFVR0RpLI0n0K/SZZ2oXrZJYxR2
6hzXxIkpOIL4hX7WrNxBRhiOgKCkSZHlhs5crfEEwNniJk91aNAPAqjMNbBlVni77jNz8rFKV0U6
gS77jLOyzmyuGJJQTK+gdPOwJ4nNfkbFrHFkDJ2a4MbCIQj2P1FDaIpNNw0i7OX4RrnaiWKxmQ3u
iF8UcYOyNkbEXRSWpqJnzo+p1AL8le0a8Hw5nqPq6ih4mBmbd+IVpM0kaqzMEPFlv+ktKeE24YTU
8p3ho8yilQi7Tx83nJexNO0hZFz/A2xflB9HRhqoRiDumS9gNgc3uMbh0CZlUK5iFxc0mo1LE+K5
K8pRUPL5PCwMZUS2NvhBhCMxYjLHObgdv8zu02+/f8q3xBMNMx+9Z8heaXaXQLL21F7jhYF6+yeD
SFWWcY/gdbJ/u9CCGN0iyeUUAlsdF98NijCUWaPdHg+3zB0ukUz/JurnTTpiPM1G2EXShZthABK5
VR450TWBjzwef5cDN/+5nXn/VUMrCusNFsOjXkk/m3oR0wvD9s9OKzZFYXk4qbFko4qZ292M9X3X
KDP8nF82xveAYJH+wCwkWATT6ynnVSgSw3t4Yz6UG7lVSKd42kG6YXmM/Dbg5zGrqON2M2IWLdLQ
NfXnsk6VC+vQqnQm8cppqS2QHiuGZ1D/j/5lBSrUgImdQr9LY4T/iEvzivZwTtYOYUHrtEK8ina8
AI8B0vd98qaMy063NdGHUrkiwXQDqTHB0PBJXKC88HUzvOsLa7YqI9SLWjW8O8ezmCTgkoS+H7al
CWNCJwXegCw3hDv4zM+7RRSLDeQmK3k/8vrVigA1z7kiYuCKjtW86E0RD9uieNm4DkIBoWqO2D32
Il29tqDW82qHTvAvA6Waat34X8EnuIN5jP6+4bee/8UHAFpnu9KlgEBo2O/F4v1exiIPGR41T8OO
We0K7irzTFMzVi80055LOsYmXtnRWNKh1/q924Y1kwmd+aFFl/tJ2rnCGtLAE/pwX1rXDvszE2eA
3QMZ+xDzT+pp5ztVw4d2hLNz5k3FHsmIvS5JAeRzQvbUNkpGTXslxNPeGFKHYNjkIdp51pFQTJrY
ncl4HIVo75bjdr4AEMFdWG+x0llf33aJlHAu5pPhY3svTNOMqVdTZ4HcnvFcBlrNaL60T9QRxuti
4ghSL2VFK6YgV+kV5Q79t0Ztx+kfqh42rbrWj3fReaI21+G15sLz2nghnfqqMMplb2c5gBvHI6OQ
qaD3wJpIYuJKQsdZaq4HrlaEAV/WhkA/j2SPNHCF+NObCz39/JLBMhyI7ycu9YP8UnABJxO7wKQz
RIRgXrfH40MblmJQYPkwDfFVwzEJ39xgGS5giA3cH/S2GNja5FLKXHlfMBEY4k1r9IaDQpavs/8G
D8QjYu+cxkYjQebXtIJgPV3rJdCuOH9FuBNrx0lSOcApBEwNqbcEbTkb8Gn+T3tfKpXzZNST6O6G
2k7SUwH5UuAEnB+IC3Xu3tcl7zdS1XSTYjkiSGJ1YPdht0OO/FerYuqqloMNsa7QJRjxGHB6Bpdx
36wFuiMudxjpkY61s7RGpF0mOigM0G7DHHIKUF55I7XvzGVN9QDUUZkTZLrGFENzeg0pNfYLOBO5
sZXPNnmZXUml8kDm9rktRU1Ku+iHP5QWqx5MpX/CrVqaMpl+3O+UOQMIrT2i+e6UseRXCdCAc6OD
qgz+Bdj1tE1TaYTMd7sWzfnHLbmOoxwVtddLiQgLs+TXhn0z4Qa2KhNwn0LwCS/0vQjiWeUVNetI
nDNKk7OPR8yrkOQfBSQEWbtkw6hx5Z/aiuvBfBw2rKEz1hWqb0RVnPwDuj0uGZlK95qulDPtmquX
pSY57h4kGngCeBgSVux4WipaCoiuCylSYIkt/mW+uaUwZzWSzimPxygHb4kK6X3Jz6lcFgvkrBfY
BCcKHpElMPKwrF4sQB3KHAXH3GTnJxGUJTG6M52GJTqzAwysmEDjMA8bGbVZLnJzJGbropNYVWJ7
efjiOsCujQspvFdALOhVNzP4/r3w0P0M6Cd2iTXtBR8+iTAix+y4DWSwr9CkTYLAllQKMLLEuiwc
NJwbj9QeGCKeOr6LIM+AsmX/ec0ieKr7d+GO/LP3sjZZZ1C99sbjsrTE5HVNRy/X0LpPAEgDTtk5
2ZnIRCfLvtGUc71J75xP3FSRDL3JofaZzlH+ypRBeOPpaPbC4PdZSal5cPq8Irrl8IlxeiPWGjXj
7/jKQKX09eb33VuEV6Jiajh+Xlt+NnowndqSfGgWypPhO1t3xQbL5qrZWsEusF1tddL4+TnTtDCC
ZRLglp/k0Ci+zBJfmndHRMqdMqS6unELao1l+LqCMRIMSZXtHyMZyc4g5wN7AoIR69olcuz74fnP
62z+AzFJn9hp+2U3VJxPba5UrXLYM66biYUE5MdvQ117p9SMyw7XkutPXmgGIdAKm8ujhJxzJYMc
D8MrtlAKBLgw3xG1Z+aG/NtEU3Kwq1jbX5fWleD/rqRo+ks2lt2/LG4Drd415bcCdio1bHjAPRio
xTSMlayG31ejLbr4M2Gr22wlAAeSq5XDBzy14yr3kPSiSUnoPsDukJkAzWXG7PPRoGBhY9u+bKEC
UbdmOqPzMqqVXj4MKpJooP2We2TidIgKBPAWfUMs7atfGRxj/AngCNqPSQAYC10AU0/P4pQMfsMH
5ZSp6jKgLb3AawKj643+UsN9fg8qtwZ4AqB9mM4rAdBW7mnxZEfjkh2+B3+7QZRI/H4mGYAbMSfw
7nD0ftJSDPuZK0a8CxeAmSDRk2iV5XOd4NcWfxZXnTe1XW68m33JeaGqarRmYDu+RjBSV7XyWcHl
waEouGtNLh6l42zV8H2zORUURCbp1sEi3zzm9i/edvIth5DaKaEAfBmQ1xZ+9/xOrX8hC5UoHpAt
j8op04qOKJ2i4hL3zJgQ20gaUbkt3urvIKRf9YEwG9iqsKRDsGF6HmexZ2/gUy3S0IThOEJm/A0t
zwaD7+TdR72krau26j/l16k7dgffWJN4mCPxijWHksifkEbE848Xab5xL+x5aE5xwXdAilnGJk3k
jvEhW5ZPtAliGq4vKMxmV4tCnByDw58+dqUU49M77UFTLc3WPVMcOiQQFbwGIetG6QezPv3t2+dC
+QP8Vlpj81kQEmQgPgnlsosx1VhNFba/l7UQJemqiKtndx0fEs/UfPhViV786+A7nKSBFzLWEK9Z
5x1zPgoSVdR/1lcgYdBhDajRqnO1OgppPHfRRWR54129Oro5rx1xX0Xjovpu7Mj5n8wzs7szRhFz
tGDUG1Cm1s1xFNkdLMfyLVGhGHbnEKnKMkHYLCvnq3vqDtzBUvqyn7re/AIHGmLWD2Qt/OnOFosQ
RSFEce2FJphtUcLIkkgcD42Q53bcLOODE63hcWDURyKdxQi4q/3qdq/TmHJxTo0VsnLDQ/AgYkwf
SkgdtmEoflI2x68yqALyxxR2406/W8YUfgw0Nfg//e4YTWKCYTCeZqG5SM/TN1BdhnwQ4J7o9URQ
57sdyyp+2VRfo77QaG/GvK9kJybsyL4OkUOwpLpO7VyDf7ESlcvb2hmhEs8ht6yK33qbJrQLW002
gJkMZ8NKP47yb8aQxyUuChJhWhPrc/PzXs6U5UaTIH9CUuuW6SEN6McnFysBeVGErxATLdtNYlkD
uqyPybfzqj2Ss4yg11ZNK9v8HCGOyRwHCOqU0OtcmNl9jz9tSA80uroX90w7Tl/nXmo+x23DpBkN
u7s26frJMiOPl6YQmTK0W7ujk/hvuymftZTC5IQi5Th+4+6QlGd9/NdmcLO1pUHkTZ4uND5vI6cg
W9zBZpNs1xJLkA3D6l0txrwv7Fqi4hsvqncvO9bGr9VKIjsaf3CoDe0dpCWoCUgCgNYMzlzjdYxC
9WsXt2muwaoUUutuKOkH9JdalrkJ79nO92w91buE0chJbE+3/KxJ96FAXziIXgjcs+qb8SWMz69Q
IYtPgEJao0FM5SwgdLIG4TOnG3+r55fUhMwtxtTHOiLz4nyvahGFjR8uPvvpgzkbC1bpZpwN0f+l
sWQtepD8e0ColhJBJf9tks353HH9Z2C9phdu5iINTI4LY14cfcsiCIfhQyMbohGX6yifX63v1Xb3
3yUlvqXz2cvqXO+JopuPjCXmrXFFOrby8eexTEbIIWqgWI0yDSY7q8ZXImIgn2e/PM2Ooc9kSr6H
XCJB3UNEZsowGBD2DVbOAFvz+U7uThRwOvu/z+maz2DuF5Z1n/kkEMVHZ2es75ahEQsCHx12uIDZ
al5K6Cnkb7Lzl4W3oBiaYtCC1ua/wELkxJv1m2oM9qdG7t7ZMtyodnEPfRqqXl0qduZDQtTstE1D
VDsJ/TCYkzr3WaVswzFawY8hHhSYIaXWshLkCaiB/giiePkEJdwD6ayBPyP3K+g3BsaOSGm/pJbw
InJm6S+HlaBc7J8+BACwV97GkW2zyPdm8GmZFGeVoDN5JDnyXDshJnhsZXkRkU7jV2dVUcbErSPX
iwuuauXJCCt3RIhcIFl951brFGLYo9p73fYCNLVi5OLWdRDhfwG1dWU45zSkOjw92qGy6ip+vcIv
BdnNvDlP/pofJ2PQoJ4X9KrbRPsUQSwTcRfyZouEi2iCkb2OaiKtI30jM6I7ctLclrSRni65Kj3Q
ZvMmfkRG+8Iz2FAgKfnrVW8+K5iJu4aj9TXsTagjSrUfj5Q8I9BGYNUF6RLS1/yCPZ28Bo47TmXv
bkWpAqkvG9EnGvFxuKGcWMS9/KZScrY4GrDbECuf8FlQf0k/8f3MOuTNhoyjwaM/uBvLqH/ZVBEY
7h+joIYzcqLU0GKc1g8pSGwaJB81SfWNOrAf2AMGLXQhGA38k8OhXuhVdu+K6/ONRrEuc31Nf6gT
OHChwwmC0Z1dimMyW48aw3ibSkc7RaqzoBmj7s5FOxuUsq8s/bItSKpOe/ZHyoRBPM1/S+i/3IcG
1faF+J7JBIgWffAyhdn33mVPNDvfAScbsUXFgO7ZbD6uyvjCeDaAYGs2pZ6ZgfDBPt8w1gkp201e
ViHYwc3+4or5LRi9X+L8MM+ciN6JYBokMLEF+jzR+LUgL1cgb6vJsmr7yICc5LPMSsW+5zi2rhuo
hrrPpDqx+o7oLfe2Dlrfb4JPJSgVmYFM29CYWTc71685YyRnqpJIctcyB8dK6NLV5AkaC3TYenLx
CBsQiX93sQlSsfbrcrZ9ejs4MRg3N+PpKylXVAoz3GpIaaB7ukcAvMPO9Kq9ZvBstIGEpPtU1LPI
xGtRqgnayGmboRukkMtOUOzlMElO8XsO7SEG37n5CP1zQKmAhLWYSy6yxS9AmljFBSiRh0jO/rji
bbBvlLtjGyM6P7ml1gGweirT9+awE32hdxGu0ERH7yVQmo8RtCIk7Kw1fPt4xh7DHXC28EVWmK8G
XHboufp0OIKrw13BczLaq3UoeeCzsOA4dXMU8qkZHVWu2rGfMIqfyuI1uaL2YIe+cl3vVRwz+GYh
czOoS1/t5uujPqbxAj+n82FgGjeg2N9MLMmC/vhgYCJD+5W7cNn6547nkCwfG0LVtyjIxQE1k3xp
IrJgtmg+RpL/CMBGVzZMKrznwaYwEcBxxXaf13S4JVHzRboghR5CWriuSPtPX+OgmE8QyS4qbY6U
DoeTK4Bfk0Rwvx7OKyOmEjI1HZEL5OfVAgkcwIeP0zM/HUZfryxj3jl6blkgOIoNtYfr5EE+Sj/Z
38GH8QyiyhvKa+3F7OSkS15yEjMJ3+ocTw9aPoCK5uFuLzzDPPRQrk6IVaP1SjvSl30y2GdTs69K
K5pcnXVwF/BcibMhMtvTHQmVFXOTvUlrTs/t5lq1BmTUGvnYyXE3Zja2NTwBYI6ww6AB1msqGGdU
OoYAP23hOv5ykbOJ+0lIPUEw9zc3mmd5Qe+bTLOYjru188hRhehyH3fRx9aj/fXM9SjICVV/H2Z8
zOj97hrr7wn+ZzkSkTBQV8Ex3ilimOHydMuAjtU3iADYSyppkAO3R2hNyyeh+PwWa7hxLGjDAGV/
1BRbf0j97k6E1C5dG+eLfa0bhhrb9ri2SF6wqrEHZBPeGR+bvT9HyKY9G0Ni3SV/YfSf25OzNQXU
0fuqnRdh9WoUi9i36TEKfVS+fldfJNDzqZxc3ConpnKeC45zvIRipybPX+8d7VosibuxCSGonS3n
fPYFiCUjwqQh6StLsLBK1EHD9LHH64fKPFCGUsUULaUJTaH9JFFuRh0DQ9TXV34vxRJNMQWl6jbw
iS6plEfAdjLYOnJhwemL5XWNjJsuVl0i5zBnLq2DBtyy8cnmvMBHJ0sppl4xJkYQBcCwtrgJpTay
XABALLE+y9Iw3LJjWIwoMTemNfdWej5CfiDspuiBHuWMMEgWTE674v85VgJK7d0EqMmaHz1y2/xN
6KiYjWSR2oVAk872nTWWa8+l2VC8RiWmQEFQwsoGyYcjpbiLhu2JNW/IGxvg+wOZ5m5F4UUt2idX
kXTuwLG01TqGrXshA1a664AMQ+LmaHrR+OCdj+EvTxlJoarIFq4VoYzIfllXUXHJ0Lq4Wes276V1
9nOgzQ9Kklaeo1ZN/LTib/vy5y/RQ+89I043xpiwpHKwB7Up3och+CLDE0XJGl6LWDFi78Y24ADB
M9yqRIPcbHyEZxNYgf9eeVwskqFwQIj2PdtNzioGZUXCqVaPGHGGLG9uAvTtLIErNUBLE/KlRlu9
0haaXXiuARPa3PwEyt7USzMdZcKRYOBK/UKQnwlYlwBOo5CUV9kKf6YI3+Uppp27wt/3uuD2hpWc
W5iHpt4T/uAFonhEegGF9SNvsm/YDFv5CqY379one9k4YolhvhC8zjAIcLB9I6a1+UbGFbH/49bs
up0Io1pe5t+4VWdxj2nifYGdqsu4wPRRUwXvyNpNjpV1Ni/hoJXkOKoElGQB1WNzgJwZiBfcJB8S
SfiAWEoir2zfjDe1tkor7CBgGQVln1gWySoyauAUxyt1QLFggnuot0NgiAWPUOwr0njJLcaJONSL
cyitLoQl9LTvOY2YIGch7JLxjyAxwpo5ceuqbuPq+kletQ6oyTp82xkoTGSV1he6PY32a0Y5bLUa
5ZZ1WIfP5aCWTRNLvv9PmWvdoZUdXAGEqxfcm1gtro7aZ0YwSEgWe+iyY03n355OWiJYwz2zJs6y
fRShBsarrq3XEW+VjWICcQgrDsZm0lSlBqcD4zjhs9Ah9vHuQsQ80kNIpWAnWTWUSBnI4mcPrsGp
6TCPj1e17ZEQXl7ylykGaQrbJF+Q7xlRkWEAOx+Db6JiFqP7Zj3c3WTbawgrITDH/noAygytAOrD
hzqENoRacY5tKklITuh1pi5CdkAvP7eeryeq/2a6gy2zCUt8j+Et4cQa/7Q+w6o+9Ri1RdD2f9JM
Z9wsGFvD6EHdHA8OipcU3z+UFOMhJDHfrQsJb5jjRYdz+SBhFyXC1CDM1PxfrEgYSQondysawcJz
frJl5rW4VNCI1NtNNtt1216L7xgOB7yOZVcUryUI2PyUA3Xo9Fr8tSwA73E95Q3nhM96n2PV14MY
N7x+qqwB4Ag7VmxdXkL44m80qJdUKHhUm2VOF7S1ff2Ct4cwtfysuCiC2LpS6adGutTQEqjL3q1i
gdm8OJ19xA65sSHkX7E3xUEBTI6piLjzokmVyAbmkzTXgNvtXbwxyu9XbB7DevcU06++Df3Mwow/
zu1ks9KKWwE9p8EhvIYAmIsgRB0gESE5nEEHU1OEJmTYRWV3e6ieElNxvs/sbqcjkMLX4+W1nAWr
A93UPXJVMax6enoUypdhDqjWX3b2L+BoVbzIEY1Y27H5xPWpcx0rmYE4pgGIXIdIe5M9sn7U44hx
xozMDiyFgh19JLSYnUDubK3BcLHz/j+P9tJxTSUeVjJNccsge/CGsirOE/p6nQoeiHCnD3W+jdGm
lr6GjlsGIOGK5VHXKq2NotYrVpUuaGsEYkEnxy9qsnN74Er09YjvW2zjO5n30HC3mxXuwSm/gJgs
7gBIjHgzooVh3dDajF2fj5NVG1TY126hA6vjJTLVDRNjGaSi5YH8DGpL8f4gY7MaIc4aUa8TNOTC
v0AogxaN7MjuWmZ2wjO51ADoePfeJoiQC+gnWIp3uD8VNEN7nPbUMS6+X+ufsui25pB4tz2CcRPL
IwMnAKrHLcxvGQpqIY+IXIG33tJKkGD3cNr9GrQdb4275QY9mNueqWY17RinlMILu+mU1tsyn7Q+
/5hVi3QRmd8UFxs91HYQOgKv4+SSWxTt3LpwtHllcmxUKMuPmwpxpqkOfvU89QoJfby7iHAKfUMs
lYSOeitZZAuomrW5uCa0CQJ4N/5Sy2pOxFcTcxkoYu+YoswhgXKD2glAmIiGNwyn2B/yO+ZJAsWg
teYUa9KRmyyKZcnsbNGjMFtJVPUTfCcctj7jsO9Rxj2qjZ3v2m8mjQy+OZJn5XyDS/5VzhyD368x
UtHy8NSCul/rqpN15AmS7eeLOozJVAI1l9ltS/gVX+ZoCV53cbPmqXUqzSMoSw1QILx5g5stu4j4
ujNDjtSKi2lmdg9j5Eq0ypj00KyDYsgE7J2XBBqFmajOEiIcPYyRg2B9JuT7ziwD38RBH5EMudeg
lcVVS2HbZ7ZBupvAqxHWBHJN/OT/KFXqvcDZtb/G62foGtaptEpsY/AQJzzpTwS5EijEoo7UtrQQ
CXi4QYOzyOwvZ/qWsfoqOiNSPKqivG6ei6PhiBrRvJwwTYIHUSttowf0gs2qqFcfOuVZVsIhR8XV
l6SZle+b9hMoRMGn1rIsYIHBBgaT1P2iQdosdVODGGiepF7pN3nxS7bGpwbDLv8YmPBFgeWwQIUQ
UidjGwzr+QO3D/rADFAItHQ0seMsTTs3zo48d3W9ss+zVPjFAzoqezgJhwQ7uu3MkBNnwX1Pcc9U
bMeWo1CY0KAZqE0FgYOkr5C3XjqmZ27wH7/i97OaAxprwltXtWUkcTnJ2YKX3aMm74vdnR/1Suol
er3Xk4n2UxsD78l27zCkKWOLd5/zAY2Imp/5qaMc0M8OQBSkHXyAy6M87faDYa+YqVMftv/mHhhe
Zmee8jGr6/cA6jNdzeJnD9TkjsUlJ8g0Ve7KofOtfl2s8JnMLlpu7AGCQu1dQBwwqXbRZa7NH4vH
UqqC7Bj/DhENwK8Pgtj6ic+8AeV7/jDSylOO5TZKTw3lSPwmQgM4vMzvKIpoJPPRdftJJmYMCCLi
XN0XqTYJ8aLrlYNnfEKU3RRPSWyjxWi6G8nNackyRSS3AvsTXIXCOiBklonT17RPSAeWnt9jrVCU
Jg3EJumhkqNuNp/LY1DvfIvYAROlReQwmD27HabrJsMY8XeUhQYdIXSL1rin0Tp4l/DAJjRhGLHz
3LVq7rf+RyhIXqRF9FJkiuKnKmsB/hTRRPbAUW8cEojGyqBPJs9/3eaJhJ8EoiM3W1swZbsJwbLN
Ta6LUVC1h51QrSoLOJxK3ARea8Nl0xhVK/Hjh2xPv61JItU+o1iUfcFFFFOVtWA5rK20jYt+t0Ji
8Grsntaesus0uhM0/wwNATyP00hD2Dgd66F/M9beJY1hxcJp27IOtyAWjtaD1Gc+DL9z9eEIigBL
OmA4fu0Uo7kUEmxuTmWCWW1Aoo2vdfDwnfkHWZsajlc8QlMqhW5KUVbOA0qrQrcIGleguiW+OQsm
uo2M0PAX/KFEdjaH2pjoq0l4SK1LgrvqM8nw9TbgUY/ZhhvEF5A8G49Go8RWlYUor6rxBcQ08t+g
QfL1IVKGkU6nNbD/Vo46TN/U/IjkOFbYY/cYyVRe4v/T3jKG2mmROrQQS2JJIEf5c26a1LJj1Q3R
G4IDr17uU81JL5EbrZIqs4LGKJ1sckorVnVlXArBgs4vHDflN27hPxNuZSOtOCX7ZNhQ4Ip3lj6I
0xI2EuE4vi+UDTnxD+hZeg0wO7l78Y6+rHm1iZSmTyn4xALJVZHH+ihEEdPqrXH2t22XUXLMgwnc
8AfKDj2brk0OWZsKn9u035ZGtKKFcsCjqqRPjgmZLwyDVwsFs8d3JjocEGjnwp7CQ+LLqFpu0Ocq
cvyvVjI2vVGP/jI01GJwUbVrf9jZ5G5ApRiEC1n9AAAQoez0iHkSXDJP1NKnRwAda8EmZ8+O42xl
FK8CfMgtNAVYwfLy0SM7E50Zc0TaY8t64vek6Ln6wn82pulWQp1Mcl+ct/tWcVeIHIdBiYbBQjX3
FYicvrYQQ3caaLrTLqksjLG6hyAqo09G2pPDv3cAsGazHdXmYKTenjQS/iZNqWrANWBzWlvUyuEn
CXMg29clXfcMFJcADgDVmzVMItj/qqXk/q54v/4PAm5YlW5tgBFhw6SHH4dKGS371RfZz418sdR3
nqPveNd6AZTFd0wc4YKtP7NAndArSdxHYqzn4/og1jUJTuvXfwieHhSnZiAYp27Gz7TN40DXyEHy
yiL+pPyc5qowcrv3Uf2y/7gsNt9LbQgzzHPjgIu2y+kdQJGEEYzoeliVQDzHUyeNA9V2Xr9p2ne8
KHl/fYg+OaVTvkS/Bk/U4gkp6ErS+c4OZ/eNRNbZTFQTvMXUltxK6bDl4hc+dkpRnKp/HkLpNfmK
+IJ4siJYAZFK9fHLLnrXoPRc1m5CDrZLqtpJnlEIT8t9Nq7PVh9WipD2EIjNDXpd5iUmV/Y2HDq2
mP5iM8YzqHEb+gMz5elg2G9wY3C3jj0R24sQFDW+vyrMbH5sgfT3ky61bYnymv7+ttExQAQ2uqmb
3WXho5xN7v0x4OU6Gxiu6afzszJO5DMzSTFegMvb4HUk59EGU59AP3yrjwJc1OfRh86GYoxQRlx+
m/J124t5/sqMCPohZ8NCsrHhqaz37D+L+Meyx1pnZfDcAGjxGGO0gIc1sx8wzZog5rdK0p9JwEUP
h66RTZ6ALfejgzm0QnSYWRP2vzAkDtviTofka+tQdFjogl/bydBNca/7o/oemdcwKvaeyE2iob+t
J4lVFGz3Cg+e8b+ZN97iWohh+m8VBkMRzskemT5XsvqFV29FQ7Cox8YX/KL+YVroThM8NKZXXLq4
ZClG9S5E0QDal/URX+3MkE0OPUmQxPUB7QFYzMBbOZEqswDsHg5IXyKWJQOR7kIbmQv2PPjeRPZS
81QeSqjkMQciZcjUuS8SxO6tn41TmaT4ptHZkMzQTSbk7GRtbhK+IhJ/yaBOKqZrTaVauuedGOK+
VMGRGMV5azfjXUdLtpJ+9CBp3AZIYnJcKSZ2RD+e9UQSu+noLyRwgnUqTeCEjXY9ZAkTghIR5x1Y
9RvFKceZUgGCkt6v/smwdCzbb8uMm4UJSXj1Y9V4yNLCKLz+5FFUmBKo+/ZioPP9WrpbdZBV3pKL
xnBLZR4bckorfYBMD8AxZucQGcWqZ9wPIDRzejgfVPOPFupKZgb/eWcKNLcMyK/42VPLNbLTr0ri
ghm88qNUdI/1e5laU5laZZHvflaOzSL7F+1VoqMmvxnQ60LDr6q2KjYCTU3V7Rkj6++v6Z9uGFol
QuDsw5AZ1YqXu3eon6N00hQElIQlo3NZ8BxClTUevxT+eaRg0ZpRidqfxRZiAmxC1msyZJXxOQMR
kiDEStHJ11lOJ53YKVpgqPIse9Ug9OYlhv6Z3lSXWUHQq51diapAr6BvcYCPBIpdSaJbGBO7+Du5
w0adw1RcTtk1FxtKRzL4IgPALsgXi43iUBPVXiHtIo/QFydDtc8ZKYrixVKKRH746vGdQMP9kNXj
N2XPntdcs2bCqDn6GcOJV0pZI+ankrVS2ngu+zlLYQtnrG3tLJwFX63nAAYiP0T7/r0jiNyd9z/G
9snevASPl8BdU2LarP3JMiPmvehYaKQV90Kul689+EUum2BzUYEEckzmv7nf5UTtTBhGMktnMqHl
mgtLkv6bBVV++Zb5y61Ev7SYj2RDlMV8x8ourRbILcJeWN8dTRLfG2eRhRpk8z3Sv4mU7mEEC5Rn
ZcAF508JxTZVTgVGOFwGcqdEanP1P/MLdrQjzT6RaERXqCU19fsxum8rrZxGejUf1MTa0EltMGtE
Stij9M2IcxU8UM6ERGEeIkJyO3XLgrSywga2unlIiRf7iIlzSQHcwms3oC1xqDtShrm/qi7/iref
utwBLWhcjFeHpz7/3Xv4T9Ck5nMtktTc/QeuVHOeSqfsDPg4aDdYbbv5DTo9qVEsPBMVS4EzHirD
bIr6DHoWudvysZ2/ElWQJn17Pcbd8OT9RH+AjOpnp8i2U8IgRlkC17NFqEWxHY/UrYRwer6zAyAm
HE4b5N37O2u45dEdpaXbu2yuSWKs0z9V8X89g4KjLeH3BAcjKCChZCFBmz6iojspwtM+K/XHPN8z
VnXU38MAih/3RTe9sVDqy05ai0xgNgI6NTXEx1efmSRJz3NHHNI7L7zJw9PC5uUuHLTzyVqiQbgI
dbJmgX9ZUh4WZWHQ25XFbDQXCv09hcu1RmW0LkWh31dDg5EcZR/O54gXYKaWlAXNKCkgBUu3LSY5
9Xn9CX/OJcl3eSdaCuCBkUEROG4jefhQ4/X/btqHf+GOmphL8lkZqixutGT7JXpJGL5i8rajrjQD
O4dIjadUep8OGmZoaM4o0hRLSRLpE3/zIpj4Qe1XB6r8CbR+MyUebjm87n0HZOscDdietgniAvMZ
AiKim/DZZ28A97CQP1KynWo8lh7/9Ado5VNJTKBlx3LnDol/fLyoRC3bt/5HbkGv9cC7eFjfGw58
/Rp24+C/Z2yqPkM8KyvC1KdNehFkqkZJLlsC7W8itUVN8TwMD4GPW+u0QQw0Z6ucob0d6cgAzth3
IPjptRdndUStIAiOySm50OMmbC7/1qm6EUjHoaWbzIu0eDqwKACw4a5NDEgU/YcN0ja0gJPBXReE
BOQPHy/nllysYasftxoVYpD048ph8SrBO3YI+YLLU0utBDwLrqJiocLqBJ7e2+t1I0HKmae7Yqj+
Z1S3k6iMUASAi6o5YKu0kHdeFVrS7y+7wxzcTzXImBNF+N9q0x9T7uKl0t/wCGz6ZN1E3icB2nqu
JnJs5mLTRMyy1A92IjfuDdUGJxouODOKpXbV9JE1RVBuCdHJwAox+7PQaSWvxFXIDeJdb966WMdH
v74mHTDb+v0iqxe1Xm9znBkhurEmiY4ZJxZauNqJGyjTp3eB75uuA13zwtr11XIoVGQt5FqPwouC
uogSywpuZchLznU2HOGIyoRMYyFOMzz1IZ5GVx1r8gdBxg2Dh45blQ/TOmUc/u9hj12iJHZI/Xgg
isDstHpf1vV6AFSsDSlJj6NcuXsuSTSmuYWtMAptF3Gx3aR71JYhJzoPDja4G38viA6MRiy4z1AR
9pjraHSAHzrkRC97GPDLvc5J3WRQ9UeiwJq0fOjh9x3cODdCddb5pypZq2KBzCAdAVKh5agMGYCG
U+80Mv3Wrsh1Xc9Pbo2iIvbkv/IM6G7IU1dB3yWt7Zzu+a8L0UD5nOZXAlg5Nkgb4mdvIEsf4FnU
BQkZBF+wOKze3AgjI+YdmZP9VpFm/f18ZfXP3uLYT3MxeaQwimWNgRDnlzkbbrOHp2zN9Akla2M1
ypYNr8LAr8hKGc+TYHBJREASkRaDVM0yL9OIayZNE3E03oL9dGX26FAW0X5Z/kIdFryfpZQplqUh
6xeR8srHxDJzhmYjR97QTebmC45ek+IRNA+sls4NBo9sgi6L2lKVQfOI/nHgbxdNXFFLQDyPoSY/
qwxGyVGkmO62n1nBiVQDJlT3fbikoXuZxgNEtzu0iT40EegHUp2sn5B6X1UXvCKTN3SbW5TEZwnx
CGbF27MvHPxu0mamj/Bf3YQ49T8CxQulvk06x0wYFPgKo2ty69j3VaYH8PHyMpoWN9mrsqlM9kwL
O6Qvc580aAfc695eGRjpS07XDG/GY5JmVWOPCIfQaJNyeol77QfDw79nKbfUZ1+cfsYxRlLi4AQB
d9Lf8NOHRJ/sGftlyH/3gJOad/pd/A5PXgyG6S4GJqrshhLVWVLDMiLnVnNO0Lf2ThWngGy5kUMB
KvP6qGu2MzQ2dIZK8VJn/LPd+UHP7EJX+Ccg10OeBLFPk2IhT4GzX5PfSru3NlOAydL5/Dh8p9+N
3I1EOz3yByQrJFsiz0dGiSxJECqQtqTJvcbGLQrxwotsm0Lb/kXy/zRbULbKZ3Rrp/aYRLWCJldl
Aw60MdtcK0GXatD1NwfpRmhEcCqiTH4LaT6e6wcRddgcIAhhcRGKsVmdEkKXb9R10Xnf0Jc0+AEb
/v45bJESPMPCENYdCvKOj+W13y52VueN5h+ih2GUPMsSTotqWyRIcbJR2rniYvQReeEeymKj0C/G
GunH9FbsNndulrcjEfnUXfyR/xsPZO14vyKmXNu9zeg6ZW3PnL3JPOFcxBhiT4SnoQznJVwuw7au
BKtsYWyOIkU94R8KfnXEwQddXJ6UQiZH8WcIb8UQV7+sA3a23KAo7niW0qTp6obBmelagQDDBYpk
F/gvG6HC5WMcJCx4C9xHTdNEJo3/RBfduUiqA4IbWvn04ESfItoLjCpJWwCKqRknmv2UXfuU2I0j
5Jdt9XUH6VVRBUfE3SM+KhzDEDAWo3s8WEXwZC8T2FlUiplgacwFo6e+s1wK8zjE14LKe/bh0XY+
XunuebMoDswX1t0u6NMMip/HRG0IpxUVVQBQz6QZysIVFZ4DFW5KOeCSQfN75GLW79zjabXPAzXZ
zY5zi/64alJbvgVDzUFuMfKZ7aT38q/syqS9Fabyv+NaraVI1F8YWK75IxdlJSlO7vMqXJTONafv
9V9deexfKbXQhg5yWqSHYt8qOzYDMga0vBviltKrErIRCQ2CLKw9bxmgPqoKxssI5rY6g8LF5lzn
a8YmCCBrzYzDoVrzh644s1hHHMUWqXWfFbknd/SbSollejC0xluddUzwL/a21qYFEYvYYxk0HtxW
7pPdZKidWO/y8vrJFYfN4xLcxhKyYQ2VmV/dKHbcdJqiSztFe4oZHKrdMh+jL/EkZwQ7icHKcIQT
pqNlG9ivG/vwN8U44pEKV8A/Zobx4jG+YpQE5NAWAFa/3UfaxUyoWqaqYmXaigU24qKPuvsImD24
QZ7tz8+H6Ci5ZjACIijxEuWLgDNnl6TxRmPhI+0r1WO9PqBxszvMl8wDznnWkdsr1Y9YfwavGXJR
t2YeHfBctSjIRXBKKxW1J3XbZJGEsvm8EIX/D/9cgPLS9cG13Kabiz5PKB+hSMh4o/hPPzfmwhn5
vlKggy1VMslsR/ito9YL7Mrn8oOm7HRu4U/kVnkIjX3oRdX88fhDRokvXX0527SA/xhS0lzMh4xi
sMHTUazXZjR4Js1Ee4QEGrnOcY4rwt27A1iMGvrSaX2o1FtCgEn5jre7o/XD/i/ITIZVMwMPeaNn
0tfaNpS6inc6zus61n0tdvk2vJRNr4dl21Thi8hA4vAGk6i59czLfmuFlfDpHen9ahCwNzl1c9Na
eLKLoia6QFETq21GI7Fq0+k6VXgwOPM+R1jU7hZeb9N+BlB/Gt8dI/B0UXdd76Ww7WhtGM4UbGRb
fl9HjQitCKHpS6SSAbU60SWODIJqAmsF3pWMA53KFMBmBRghYePZgsKYxQCA+052JDBbgu3aetMj
KyzVs6ZjrPC3g+8ukFKU3dffVzCFpLRsPSNRrsO2df8hHsuW1tUL1qELFjzIfPOesFtOI4erroYj
N2umswj7tCsTXljcGcHVK3fU6NiFWzUS7koAGkRq+94iaTzNNQe2ueyEqANDDdL0Vn/MnBrvhlE6
wMTllRheha+u5AdGScS9AEBaQrsIdVf9r7ky26funhxhYIJRUCQDrpcZixw4mdJRcq6QpJlJF7xv
NiCNV9fMLmHpdfVrZcAL2GFm3v0u6sg0H3emlVS/HxHxw8QuAspa9jfORUdjgZdtlyaWUPG8YBTn
3IJ+ZRsXQJAOKEKvMlZo5xxyV0iqXJbiU3oopwpnHoOnLpjQgf3wU/PmlEvw1AlUbKnrlo0Q0cg1
cI8jpenxY79rM8RvCtVAeu9Co65W6HfCCo2fY2yYLdn+uhJXsaepYMUFhZgLoQBEiBcS4E8+5IEG
ZFnSTi/fWtZtAXv+U1jr0oNvOKe3HvvZluyYUZjA3TeJEFgr5VtObaB5KRSUsj3SRW1bALCXldKu
68GHQ5R4q1zzBqiI/RMLePqPKW2aGymikjePY62l34shUwF8GlD9df/NNkphifNKreR4xgMxHPDI
IJpUv31mPTCgaVWulZNGqYIclCLQjnqNHqV9wkGtESwBohDomImXhx5H5oTKwqhKA9QuDITP5OpM
beqJ7OLJMWhDSbO991RrCQjLnqtVcZCthKuykUoQGAmkjheKT3EEs8gBIVFac0DXjgXZF9vs6kyx
/OkFXTFqhFkEl5STd1lnPNMhELKKWH1fch/blVNOvIDTi0Uk3XAzBri2JOAvZ7N8fzfMebU1NaUY
mzzMgCdRHUo6Uc3VXafL/llbLh8A7KpXPAe62RnN36E5OUENEZhY3S85z6ehKjg38Y0f3ffzN6uN
Ldshv3RmchfATFe+hQpuT/niYGdGvmJXJUZunVp9GffYaOU8my2zJtBlQCMRxvYSSdK0iJN83te2
8tqW+WYV2yc0S59Cee+m7oDeFvuSJ69j5/Qz1gRsbmoTERS51R5I+z4HGAmZ04R9zZp6rV8q3Vt9
vNyqLg+WOJQJxfp5STP13vdg7kyt4RFbtSffb9vNbYYSjY4qBNvXlbv/NSH3hWceM+CcB0SXEsmR
9tiDBZ5h8hfGKL0OPhSm0mO3Tib1csGz1QQTgOS9v3A1/AjZE657rw9qP2Njs82lGkNzp3mMNPQO
tULgTmJcn0kOyoCTPtDrSexpUzD0Jp+gWffDtv4Ps3obyWwoVT+qZ75sz12JpLDWKAi1yspxUBhD
BgnKFT8VgPp2EXxccd6b7FUl1tMpXrlngPR1pSWM0jl3eNgNSb0k8WlaFsXzbj+5gYd9d4evFb2q
0yGEyK2q0t0oazgmD6lurROg4b6Rt/RkVyumAwsTElFWZHnic9f7fGkIfOYUWfZYE3lqI0yrfAVv
N84p9TwNa5DTUUlWKUMSNaMB15h7UX8z0QKyBiuQu1CdQ3tuatEypdFTtTFKtCnCIulvDjrJCsXo
uB5xvw5wXEgjzViEHO3XHopnTiyal94wglLNAq4R5qU69fk9qEpzgWxXHArEd6gdb3Y0BmClFZPf
9RbS/lqwARaeLaNeWxaLV9Bv1XvJG0wezSpOiLwdiv9GBpOjO7nQKjgBiNrcpHcWNcYFLpUCzS7t
x48a37Tlx+LLnXejoHMcljrcSaXMx5vcGSgXuDX5hXYhEla5Sa8Ks40QDIyxcAXySvfpf6/Cts+p
4aWhvIpx83Utt/Oj7quYUWT4f6EDoiVLOuoA/ACnbxehHEXVjrNfcdcZ27ifH28lyUN4CvGiBh7V
oF3sZIiYEtVwS82wxtGciUmec64i2hx9Oo0Sfd98D8yHZJ76y82y5U4nBpg3YRG1QfaFhZPqpxMJ
tZgxrsKfyy7kjc6bhAHK97MX445ZwMlDJcU9Qn2uf0oHIwWdcg/RtywgzzhuiTdwI2EQPWr1+ur3
gr/NqD7fqEtYgnktWOFwuOUg9aEPj3CmnHeX042WD8/IMEFxoBcpCIJ5zN6Rttoqhhn8sa7AkFiK
Ff8uut20V7PM3STmrci8yRxeqZq6FkfIALLesziM7MNzdAZ6Dh2LxcvlpZgqXtxqiu2LcavU2yWj
weacg/QaOiMga+hTapgK52gpDi3UlZb2xBWx+2/6S7Mgig2LbN0PfZBoJaWLA4sx6ZzYP/GEGJJ9
ibNKNyl2YplNdzIgmyjiz4rOzHPVOeMmsjruhIuemXyQmWDAzu3+qkD/9e1Af5WIol5dmXhNCk3X
IXtZICaek1h51LHQ8R+T99qFY5XPll/3TAIIehcykqHmVlafIyK/gqElCUqJt6eiKqfStZVky2L6
9+FMAln2ANlNcfpYq8AhBYdsqwg0VD8eCiqczVE99+N6dCWetzDix7WlPakwKhBP22qRy3vUqXiw
G2DXZMDlQGciZsLfYFUrSY8jetSJTlFgpXnl0V8AdxWCxh49I8ScdAr4BYvfAXGeL8/wLckPApI7
1M5MbmvMvxt5W9iwWT5nQjIO7g6AXsMwjYvFlQ2HNHgd0r183pW4n6Mch6j5pu51tGVPAOX//Jar
opZ+v+i5yEs2Ne9KwLmpaSb726EQANODJUx/qOui+z4GgEDWrXt6Ps/PZEpsAF61bpvtx9akI5B3
q9XHG1RL8dkJZW2oDUVzpo/sA7/qmwaEAnt+gr6xaggkA7IDpzCy239QaYrJN3FWnjJ4rMDd7c+u
WaHHGh3XSQ7zI/X1ySr+p8Nr4EnR+2/Q8aT4TXtU6jZOcjLQVk3Hr1O1RM3Nb05k65uLwPWRH1mh
ADd0a1UPhxa6iq2O/D54jjKL6u9mAHpnWASM51GALWZKG9c2EmltaTLKJy51wXhJRL5YqEXpjagN
XSSBQJb54NSnrvhB6CppGP8P6NdBSEsPYCQMen52SLjxCQxW5oT6J7FkMXaNTEhgqgm21f9fzx5O
zFszRjZ4e61E4ewF8XBZBTKWG1NvUlUV5QlUaPNJSgXtTmTCmYB6I0b2QlTvxOCuPsybkpu/gBZh
IbwC1ROq1X5DXe8F5jrjAkd4jPwMxuv/prFFoivEKGhgfOs9GkkePFSXqjsrpY5kfTFVxIlmyEoF
uN4QOZvbpcWtAOPoJNuCrYRLznc6jAutD7QVOJPImIWJKhcxUP1Brgne946rZhFvaESzz2BGr9+G
LlNu8zw3RSMeImLsERGqk8tDjcZNQzrfmxkgxec29PNCB40rLEd9/pcZqNoqVJd63L7+JIduz2Tv
rABwHSdXs2mPGBVd5EIWEqeXcLleE62lyEABoMkgQ9C/cumZZye78JuOi41KHrSJPGSLmiQi+dS+
PIJxGBrlpOLiu6mL1qSrxcWtOdBCsXvGveCTofthY2HPqQWclMhJ/qOciYTeY6eQMIVlQVTIftDK
epnjEciuaTSAfrzc1Xjn3xzLru1TpAes1qvRIapTN/xClHo5OeAQBnwkD4055Hk0kaES0VTnxRzC
G1yoylLQJkayvxPalq7uyEasxOu+KWgy5z+GZjrMrgwe853PQd5MFS6b2CcBXaXkOWQDzcgsFYUf
X5ZKDdqxxNaE0ySjfGQ77frdrCNOdIdum687WH4LLVidqrFDjTI8bctjKTGXfETo4VBws7oLEFtb
aLH1fCr39A+ypJlv4keRi+3qX3PCg+/vw8VjyH99oEfepafKUCjq66hoHC9AlZ8Tsmp5AiqqeunK
XaqXoV3TiWiTmCBjZyXt4f4xuXtgKpE9OyGTWixNRdbsh4kFjdJ1bbklkN1zJNdJGmyYgIEUp48K
rD/DL2PVdz4NcIH+8gszwjgbnhTrKpgVssATEWl+GzfXxZLLy2Ii/pDWq3jT8X4C4BFBXM54WeHS
xIWyvZquIKUDrbJ/0utRP+UiT1yrzDApph2v8XxnshTi00wInjKLYA4SToILMDVamrAg5BuXKgg8
K4uLuN1NakOSCfxlRL7zql1FB44IA7110cpB9yFNEmrqMWcQiVSGNWughQWb7+brN9wgfxDJrTOV
QSyQfa2wGhh5nhG3RIcGAkQHc1FqPT5F5ig5Pc/LCKqrx8wwJu7v8KRaorBtXsBxYfEJgnqAo3KP
ferjcokEQ4thVLNVF6KyesdcIJxSFF8ap64CDlNLyu7cGateOLxoTaIZJeUyZWcItYHIP/guYRSR
x7D8q4hOxiotlEIHUyGBGRIAL+AVsaRSmsqm8ZiSNmleOYTke9CM/ivns2Winq2+A+c01odT6GTQ
mGXIeiNT4Y8oF2pFVmhNQMJonaEcLcP+vayQzBvhB2X6t6g0+GQ57IggCAx4aWFHvHXngZgUW3Oh
M0Pn5JfMelgbnysy+Q9wd9L5fFCecMmhIieZMEFEUh/su6Taiv5s22qwAV/Frbd0YzKASoZd7mob
7vXMk6+jNOIEBg2eSjbYl1W9/48fA0WZsMQZ1Piswmom4IuuxB0FwTA2xbeG+9rVjgvO0eU5Nw7D
OG1n5Fu2MSziXZG2+YMxQ4KkPoehC9CMqvWRhbd2Pm5Ten6uGWSJSMFb7UEyUTU4vHxa8qvEcPrx
iwP3JKG+bIZcLjMGxeH89lwLs1B8uvW0fCtg4kM9fUUzhpjynE6MMzRTR4CEWjCoVvQYQFDRYZHh
dkaiKfIJ96w0Iz1Y6BEPAq9K2okKGrFy8HIqi7mxFajNvNu4EupwpEO5EWbwSNjFYnW+TRMP/RV4
Nm7OagufdNsIdiY6uymrHBmczbo7Ls1ibBnKyFQIb7JNN7UXOy4OlhKgwkLkrp7j06qvf+C1pNWQ
5wImgTehWHAI4i81ao/PVUlXmqqzuJT/I0jWzuxXeORYojHTV/wBOzdMdvCzEauD2SK8M6TUIxpO
KI/0GUUQR3ilgn0VvbOl9RMRhjuBV/Cpii0tYorNCNFJgfy//aPicVx8r8BWCEBkxzhVHZuuV0NB
rw2Yo5ehLWWlKbyndjdgOeGV6/oydLINYo+A7BQGWPzHzW57Ia329JMv+IxcFa/SccWwVAP+GTkm
i5XMvOy9n5psx04deBu484Yw6hZPLmy+BMjnQpxlNmxudUkQZ4vg3H7nHqOORsKIwR8xkFbHn6JK
koXKp/MyPHfi+F1re8pWh0X7Vt40YCOeNd6LrJLSzvfGtFuLqEXLhCx58kvjzhSyjeGXaY5kX9jy
8zMLsLpHH/u73ogJtp4umqu0qgkZ4bNJyQ57fozxTlf0caLAYTz7gyFpJ45VmXy2ITSc/ImaOSFF
55bm1HFtcJUs3LAO94JsGDCHLuKaCzV651sG24N923PzAZS4RnH/lEDepYb6OY1Vt59AOC7Iszbh
W/ZZPh/hme/G832SW9uIg2hoGsQtVuEhbpzVm6E19XzZw+gcdmyoi4+RWX881rWhBgj/9skB53na
fOegqgubboodIWxcAYkJ98NaNzPR9fBTGlHwcT4AaJPZr1b4oF2Fsf5eacrG26nUtLIFLoNdwcSQ
zC8qY9zRc7niH5tu3cKEfe87xl/dzuH6GHxvs8pcKNWOhu/+BOwuaFCnuV51i7UYjeWuTsWRsVar
2vB9l6U1e0eTh6e3oaneRt41vBQYPNIcaLSHm299pdnOae73FPXu45I98+lZ52KqxD8CBnm+SG69
JXFaNAo+FVzDFzYd+QWfcqaDhgWTLp6EC1ZKeLNis5jPVoHRadUzpzD+A840zi2uzA2L/co0MbnI
K2tPVkGxtHzJQATcxNguxwDDZEwDoGMZsbTECaULfagNzuUG88eom/rjZ1rGRtylLEx0lgEn9ziE
3sqJ7Ri0QblL038NXr7fHdRHcEKAqnDT/Glm61ktzz3b3i0x7/DeS0HO75OL5ZxoS1lsCQUI4LDX
ru9pO7BfF87SfDVPb0A0fuqHwLZX8cZ64M/NlV8bhLOVxnd9kIeV8kNDZ7UkUWs/hL0yMdrUcmki
PZhqZW4rtSdDBl5xFhcwT7YI8wxP9OK/XLXoCqQjRULAVAv0gSOcpBcd/8FrHVnH9UxxHR8bYnto
cC7UwfLap7NxrTKUTF5aR32Oj6jklnPZVBbJ3IuxOribru4fZGjr8AmPj/CXOLbxebYqjawz1g5M
PXMHFspK9tiSaoubUz8ZMlFS5GiyV/GRMk9d7WDbu/UI0gsiZnBfVSZh972vnIZSfOFpiHCIQLZe
AsdgOI5HHZHYAD6v38LvTBR68+GQrz9QhUIizZmdDdJ0nDPsZKZHbgTJVKws2ws29mwIcSkW4CPr
1oKTgww0RBz+C5minK2voIBSVJdjAmqhuLKInVrVB7U8INC1zSDzPRf6XBYiw3oWoes9U2W0kYJa
5Dc1hCghzdyagY4EIDOZNYsmowHoyAkOzv+647ZV8JnAI9UxWt19CbTVGn764XeMAGC/T02SP6xy
1bh9Yfv0Lu+LK0yBYKFeXmNQQYehMpVmjcrYTL6Abej92nYxF20wMToZ2Kru5pchE+3zR1JW8HlW
+I9/mZfzg/lR/Pe1ZRrg0VNmk2+7G413jr18XhtUP+PZXYrZBDDH+TWnLNnG2Ovgoa4K4IXI6E5+
NbuZWewfbavvT87V8fHarcLXUhSPZkD73VAN+QiNXJWIra4Yyu6c7oqtQ/66fjqYvjF2auTAC4V5
RU2mXgDuIr56L4lnw0MenGFRp5dcdtAJ+twCIavTrjZyDtjkfmalXQ8TI0v5PfVmJ+tdNGZ4rvHt
mXVI6VDezfkHRTUStOQ6665jmHATSLasAZyx8svrvdlnhTJya9zP32zKKN3ftQsQ0PvjEmYEx09D
5Ugpauv5ex+X1evWcSM8k5u6adoYQqTmbvwTq1I4hmclku1rfn4L3++Yan8iQKUPuZ7teS7TL8o2
TXdzN7CELduIo0kqWrxkXfbeoMq7oJdyj54Y2lx9GWNitf9Yp3bR8Iw+1m/sWyNE28rF70lCh32U
gVDzWJ9qFVHsbH7fyEFPG29mU+Ia4moyr7XkfMnLHvHjak9t1NKPwgC4L13fKH8BrR2DnrlvurUB
j9V6Py31RIIzqw1d3UD8lGN2zARpsvrmHRu5j9moUbDZ8JUJqz3oa7hx+0eJlYNv+PicrTuaYQjy
N2Id1PqAsKjCybzpzoZQh/5eyTCAGmpBwRJxiqmaTQvEgN1V7XxHtZwHIMs+YROumawf1e6+CgBQ
0GdNI5FBH4WqH6Bgy67T5pxHfpMms9EEmpv1xLM7kK3+aJH8CN1RbSXFf3dd616rHhyT1+Ceoha4
00TjGQCnLNWWdGyH1NwZ2bfiQgk5TbZ2eIoCogpXXVr3QCyCFgsde8C3R/qYgL/3FmyJgR0bAS50
Cft8t7evdJ3FY9TerYqiX8j6N/mROhbhAWrAySjh7kRKIwMj+uPKfNZgMS93uz//ODr+XMvyOvXK
kNBtlcTq+f/msfi6s0Syiv/dqSPWDhgWawkPJOek0NYWoTpRJqzmGuKcT/BbTbH4MkqW5yWsFOjT
U9i2MhUUUC55Ju0dIAs6/6nPCMWAlvpKUeZdy1iY1H8ftqXww21y3PaKNdeFpXZRyzio7fxtnqKG
s54UCxpOtD+6xgmFp2Q4brqfWDjeUNfuWvaz/WAmvFf/giR/DozciG1Gw4YBEzLzr54uzbrrut8y
XktAEw3lhNrzZ3J5RW0hQha/rqfRE0HIcqbo1o8gPwwlX5c/sIiaX4VcH06+jeN2KUIgGcIdT4iI
EKCX2WJLO4KuuTYWJNVzzEJIii40qptPEpiAFZGKbl53FvCzFSvZxEuaFeI1/6GDsBrbOPaw5K/Q
V8XaJvuGvYQLQ2X9MHe/L+W+pC22Hp4dNmONj53qUVT1q8eZck2IuYKGjaK5O2GwfdRLslCs1kZz
5k75ZRfy2FAt2alX/RFiqWXCRHvFpwkBNbzcAm6h684F3ZTxu7Fnh8FTdfAHrz5DNR5Pu7YkOJP/
LKZU5eyeWzNqMQdiX+TNowUQVuB4Ce+q7UdO4FAlKoVjbiWfZCEZIbYxsQ0htkdH1q1jI075B8XM
Cp1ldj+7DDb663k9zv9Qd5drg5hqUXHX+0Ps0/XjVYPNRQbEtaNslmA02B2PV+HGQimljNdpnN+q
NVAIAsFjunzJgfuW+YXkBU529ws8hj+oFmZR17WzKi1gX/1Q0SHWUmRreLIABGZv9DupgfPvu7ZZ
dO7t0290KM1OwiEoirxALcyNNpE/KrpqrH5yix/uOj4946y7XwMQaXQPyC48qFW8T7r2ro0sp5oO
B/lRjeUSy+PGVMSU1D3UhMJXE1sN96mNzGRhnKWeyOeN0cdw2stnansISO8j9i64jTsaolat19es
yNW3lu2HCvvg/lrjTYrrWua9Qzb+7SXYm42U6I/cf2vTKnqzLm4P3Vd5jPtR+iD9nHVrIvhi4/37
1KWr/Wf1mIUNrz8gmgD4gxaxgmCE46ZQLY2R74lUdWxGKvg74zAR6QW4VRUHYQlPlEtCPotGE1U7
Mz83Nlym+6VHdhBbJ8M2MkWXo8SRZPWU216ZK1A1T7A8COR2g0UOZuxUobwXhMHwTXGje7iOwuAJ
PiiaxhkT223qHzu1RIKozItlgpQeoSMptK5BQbecY7KLeI45sCJDkrqfIG7AJVcdShQYkS/cJQkR
WCL4lMjQ/8LAJQwUlLLN6z/d/IHyJ4xVdFUz1I7Nqw5evmY+H6eq/s5KwfUkGSteYREXi4z0lu0m
wJctV7usm0K0RplPjhGSa+G1wMTRnKKeydDygRltdjhCjh1WJ81Rg356dXcZXnIMqj6Zmeof1xkS
X4iXtzlnoOYK04kgVPsgbouH0wNDOF6y8BaEvnyOjJAXJz9HTfJP7lWkwgdSdSxoI+AH6trkTG46
YJ4EobFaulfbo7qM4QIizHt+XifJvGFx2VmwAk62SobC6TouTNI7xTIiyO9RbI9bYjvqTlbNT2MU
y8JQ4XiiZTvkR4BRzMxqkLjcqsXBs5H4C0tsLsM1E7ERb7dyyCMmS781BDyreuE0lnP3Hd6g56C4
wpz/hCdpVso75goy0Gsm4nlFVcxEZQRj94zg6ihgIxghVolxIcFCB29oPHMehySl4uXufUP0tBXG
8nkjdAQCO/NynhSgoOwa5KwqW7OV2Bb41yUdVivfhxVizs9yWRIzMsHCCyLmJ5rVnJVeAmrIIVDp
sbyJ+w81uhRfnyVrzj0MAEBk6fWn2I7UOJgWscz1Qs5TCGuJ0xYQsbuxLjJ36VWzhXDUz64M2L9H
9uTGb9Fy+wUEZF8+Lwk+sq7+LUqf2paju2SIvB9HtwLDp5j7pdd2U3g7l5/XmmHGGim3uci3IenV
rp/3y8fOhFtt6d69apaAhqoDYYwbD3ngIy2qVQZPDd4hS4MFVBwKJO4sb5TLLgnRS4X1r3E4VoE8
ZgKdWMCGryDwiz05qkyOYcw6/Y0hMYT9nIKLCMXdyNcFWqkuWpM1A8sE9v7nAW2KkOviN3eiTNih
q9Xb7pHVsAbh6twXREGAOwELzybhzfIG38yZyIvgcQhweVeMmExh4SnwE1KRyHKMBn6j06dMl06t
xykvLBwbPHrUs19FOM6ukH02gt6zp1vLW7IQOhXNKBDlRVdCWVV9uFe26STCIQN5dHGiV8Dn/BnE
vaFjJlxO2vjzYuLHgM3xoHd8YUaS/6d7c8vv+blloWL/e1UjTpd9p2SFoMgt1Bqu6QHHfzrRIJog
X2LMvQgnjTnqpCge47JH99gkkzCH6prGYimmWYfa01W6mnIpNc+bSUBHB4aMObU8OdmfgAYpi7jb
rEVK88QSq8x/JEP8MiOtzZ0g++C0IK3aq53fDv54vqEre6/ei9/GUYdap3IA9/4WG3tTvZfW02FQ
4TRFXXxCp8cD1YZ++QMVfUrzdmytFjEyRgnzBgRVroo7VSUSir54QqIRzyTVCkxfItTCPqVmFojr
tDetQk0hMH0nT56oqq/p1yOSeJAD1D4aDJjEuOQDkwDGVLr1UBYAD5XCsp9uoTKnzFOQl6bVnCbv
tZqYw4etlGOC9S7PxIfUNMMe2ii7xmSNCJVMWi5Yc3mMHsUuHj2VYvhturU61c4btsLJgosqX86x
m8Rf8jMz4Qi2BiKRYR3qT3EwDQ8i7NzFXUPWcKixElzAi5qi0wIZmhgWZQ/bqDHRsegffwP80Al0
G731+vg0TYDCURG5RSspP9BKn7GUxuOE/IDPMrqDAgTVM6rIyMiutpL6XTB5d0/B0NlW+jT0bT1L
QfNg5P1KUZM5PSImPdAnbujrM1EL3iXEvGewfD2GPgPWhS/fX+WHAa2Hng/tre5EytXoEDwk+4YN
AIXuVHcsNW7WovOhK3kW+S2VkoU89/R5Z8jZSc2L0x9V+JvnBU1/mZ/Q40Zi5LCPA3gAa4eMkLG4
7occP8G0S3udoHknLHOgEjQmU/43qRYgsrGXXqMhiZDuET1P5UN9ouxODB0GHx3uAep4ZNymdT2B
x4PhSv6YnshY+tWcB3IOdXPHziLOM9OmQC4SKDJU1huz/9WQcHYbdKVKR8TjARA9aoSppRgapAjV
opi64Mo6tCMWdyrU6+m8LLE+8FpT1GDkZA1fOcZyQT08iOqhfttEWAtwAWym5RON28cLbHSJf3iT
tqZ34fx3QhuEHwviIMSKN43WTQlOAJidsXCumJE0WL7iHG7dcYnAK8Faab+/pr4VoPA/WCfwEsP/
C3D2x+TwNbmQV5h+NwgOoZrvwz/W0FKBtEMSjINQa2SQ3KL3a5m61RprkVtnn80vXIiOVoM8G8z2
VhFvJb21+xFZ75Ioimh/wirIZC8lm3fp3/O5eHA9IIDqk1wDlahN/2bdwwUrnhmlx+UmSAcorUZa
/B/5uRfvjw89Jpah/LL+0/t5e+I3h6VYBhm5Xk1B6Nh+MRl4Pzub0m124LHp5RpXSYicBMJTGcL1
uoViLp7z0EPqsciv4OtCCgzvKZFbsRzLGVdDdFDTaYXCllPze3telIXsPWs9kcjF5/kM3zKoaLeg
1c1PNCfwhUMLFbSCYEoI8FkYE4SiPyiChmNYz0iSlmiVcjLfW52rYJspS9MRfR95DOGab9keRqIV
NSD8nGhMeuruJFcVwIpNy8c269xi+l5TLEPeVwr5Cuo7NNoIsiDn0Smqhr373UqptGoI/dsbSueu
fz4e9Z4pFhcoYih6+270S44n0+gnvQIRswuBWn4Z9Kwdx4Fyxjavm/kXUrD5PkokVDmlEqpP/xiU
KliQn23i7Gqplut0WqyEpUZLxjYB4WOAoE1jr8A/VoKZK8uNso8xtltaaN8gCS2ekclni7uMtQh7
4O+/Ta7ANV2gDbuIRlGfti7egMJwsYrH9GpuK4G12YlJmw/vZQjDK5rPn38Gu72tMwc1Y6Kvza3j
uOrcxXkIs0g3GNgdCjMoweB7kswbeZ4qIfhjOm6fr2MFJr6wVs8Gge7uazc4e8+lxUvpunU0z5RL
3Ax/rxiHTy5dIGeTLt5gvLrznfjQTxWiacPUF6csXYFRlqkiCmCo++R09tLfZ7TVjKujb59bCNzT
vImv6imoEpjI51BlUQvpm965BEkXPZDt4RpMUvH1Sunf/1Ysyeuaqsg6qd3LzrpBpGrW70OdAaqg
JcRRWVXUwuTVsqo1/B/ODolwrXsqPXegyCp/YGrr9GHD4VPpLGOO3hrChKEB5u2QiZuMzX9abt4l
6+ttCE+mhcOyCPrr4GxIDZYIhtsKMgplPUfTxqqnZJ/jjVTI9P0VfBdJrWhdpwjRKFTBx4N5thiN
MStGThJT3x3n11RUsAnGsS1NpeMpxe3CZbxqNoS444txellx0PJ1v/Cu4fOEHA8XQjLuzOfPJzub
EfiDctUXzfjQNv19NjdXVZkRrqO3HS9JXFlkkxhcwctkKnd9ttMMVY4AdbpPXfVdgyc6ihzDydZx
1VKhmbSjhYwJTLsv4IYQBEckDeWCXvTPQt3P2yHOa/BDT4ZsEPB3zFixD2KNw0r8ASteLCYKQ0aj
H6eEX2YrP66Qqn784Fe6it+mS53w+AVgK432xLSPOC/SJbXIkqjn73EDdHSxX7yk1GLs80PuYzq8
ZRMz6OuhcLJ1rZQCuJzpYlmZ1MkA9YpyM+DkN/T0l8/lVh0vhdVc4T4isqx7h4sXM3A6rG/gH7o9
xRDAYIXVa5V1pGVTlzLxWIxlTQ+5GmSkP90f8Q81UoSH7x3+T6rnIRwrSDMH6Wc/BpDpaq5KMrLJ
+QpYQQZsDWMM+5WWDODTdVrDbn1/rUBTFtLSz4k9QfYmA/HEP8OGAoeWQwQKF+bVq0QIEKYat6Hc
5V8GWXJLsKL8i3mXGyZDVmnPZlFb2N1F1CmqiDhlcW/3azG9+7hrSny8IgylL4OCft196qSha7Ax
+ErrQcPuefL8ufjHycg2xHKfsPahF8moxvRzztBj3RESoyG4RWKRug/8uEo8Y7jYAGZS0Gr6dqK6
IOlifwGD/s9TxN08Lk7ERaR13HQvh3IxkwRkHbiZ4M770YIz+m3OXXtOeFZLxD0Z1oqo8JmQRVOn
yFAtXZU+tH1ApXOljy9htvpsM0MHX6ABtw9iGi4BMlRnqXE6ZJNBZUzpb4Dbpaoco8EnWqZG6SaW
/l1RQNjmNMensGtx6zfYAdCW6HfrIGLm6do78B2CXdBroTcxgiwINvGVG1cNsJ41yIU78CG6bYlv
coQ03CJfhcbIUmU75Yu9Gngarlf8FaNidoZWSTn7lpjAwo2+z0SX79wGWdArQKopomzB06OASHry
+WTI3dpS4cQijQ7mROovZx1VptnJ1o/YzeLdcBZfDR2ykIF80jj2jiWRKas0gTKRWMIjG8hVvSQ0
ixuvpc+gkipOGCbnUVUqq5Pbh4BphhdJYXtQeevdNoIRoOSjnSLWY5nZaU3OfhKFQ/ctjvFMYvhd
j2Wev2VkKrd+k920aRBpAZj9T7KVLlGi8nT3h/fo54sCS8xiedJlg0WqaCBo46wF1jwvbuVdFdEF
7AhiJW2ohedrnMyWitisDxalifAECYn+uvKyoXVj4tpYRYfc5cijP7wEK90g2GNFPoIaX+L7BshW
arY/S76KBkOHes/RQbwIRIT0VgmWdzU3QRDVbwDS4JA9HqteOtD0IQIrrakyX80dENXmdEZ+MmSV
A8d3KBLK507NWQVHlryQ+q6r5aON1kV6QdjqSyc9OxrLaxVUVdv1K1bGOv81Kpb3HkRn5Hqjnegr
kiMSw+p+4ES1r/gdUU7Plg2ZeOUTnBDBZBOIcwDWbdDnKdx/3qwUtvf5qaCIyPtn64RPpNaHGuuz
XP4IXFBTORRfNVDVfl5I9PLIcQ8c84UmMyXVQK5TOz4codTx0w4xTclVIQJ3CFZJLkjB34v6Ka0e
snHyJSoLZmEOyaa13R8gFzaDcsDWtlyCxdFfSBrgslH8EiyWezT/kqIuMg6qGJuzY4P2oLRsF06n
ijBe99aAoEQMJe7wLflE3k/w1otTmi3/8XsmsZcOMkrrTIjXf4TVm0kWL1ii36F22opZJ4wqbkLm
m8YpUXClrwMiKa/wsGmZhdm9GODZJQXLbcd9q/wLPe1bB4D+hLTkBmxWGntIuY8raeHlr50P2zv4
8MfPc0OAP5dOd74mvhhtL3rlit6lYKVqJqpA9S+hsS9ZlwlNRJHIPAxYNDDjOL1fMp5SSa1QBJqc
mJESJ4FLwkQsEw3zgouN6gJlHqjDAtg82/vf93HAVk7Kxa+rmz38Elcaf9PC7x6XoRUvxQdfWHca
XPTJGaIjUt9hsVQ3C2NYLS35SBTKEog3dFx9eHTmQ3qD57YlZMuDmRachjhV/w4QVMi3En5UbdYZ
wZeOFfuDIhFaBhJdF/0qT/ntiE1Zi7cUGX8Jaa1BZ6XLr69jHR2BiYTgmuqQjMwUOvovo0AJJacL
ozt/cuGT6Y06fxW+TmphjylP5v/OksNfFHUoXm7nevYAzHX1iYK3TWiR0qgUP/qyPsKB4i5KRqxX
qIqfo2WiFk+w0pBCDdsNpgXGaqmL2dJMv8LEamECqc6l/rpL085FG35degs+Wwk3nBwWoagumPfp
LxRkpaFBBMsfun8cVQguvTaCYO9vCnGLvS6k6ELT9ehzQGDQ4Poa6N4qB4HNubmvLTPWFWr9olsW
zeROv5seYpnyR1+Igd7bjq685RwtjjGaBDvA6EJ1IL8N/rdpbzHJcDtF/6kk8wBEF5HqBNROHqTk
PVEbUJHT9Fkw12cPn/O//37aUDNVMogaByd4VaydXE/PVdFNEMdL9/70nFIZMxGWNJRicTRxdgvT
eiJI3aBw1bzZE7mTenKdEnGwxsCh0XLWzj3dGjZynnhmkR5B3rac1ympjIRjnzlWOWDxKspDuRFC
QlmK9ZLJSyOOJATTmxsEgxvQfn9r9+6xE61CLcnpCn5kdKHc2uaQ4L/Ln1LlOhPQMAvVuRUq4FbL
0IkYmh6Ewo06buC8Z5OJiXBzGbgpdllHCfhkvgLUWY2DwpD+4BM4xcjDsbRsaUG/ph2xCsi0Tfbc
CFdNs04eChbC+4s3jA7K24JQ5KxU+kTd9prAw8xR6N+xv64mMytZaXq/DtRdd/ZL16RRbDsrymt1
L5k3qMC2w3ItJ0I7/hYC6oZwUdLY5jjEbwE07Qeq/YSZwrOKXwzFmrqXUbSJbQ0zZWKrEu+y3T3q
i3puYL0spbt4UnP+GYHKxCMIPXn+cYtEunkz4LgViuVGmqN6aiq0xGpS7sfn75gZnqyE2ERgFXYk
RcTByLn56Pmu7ZSTRZa29TtNbCsV+qgL+n20jVLv6uPc+Pir+IiiO/Guhzkg0ahp5ETxBuayrAjJ
8e8fjUCXRgdtwebJSQDN3GlgUs+UIVGq0xXAqGS2MaNZQD7xmJEENNZ4Gay7yt4oBhnd4MTS4gc3
69t3f5sOoPR48R881WwQ1ticjAUUR2XHj/Sn622A85fzeFkeBnkfJ03ag+2PGvmEWkk76DkwMt7V
E6NonD4+rcXHl8tMg6ksKnIle4tgghnwIl8AXuepBsl6YHlZ/tSjKnQI3l+0wTALwARB2i0mIZog
MBIeGcxJUCZkgWmHKcwgv9r3GfM41WMEHL29GiI48XOUDFjBNVEmDEE7cRWuMzBThQ+Yr4XRqEqo
lVBTqB5NKCp4OtFMsICUHzGF5+dtoUxWgAfQgYWgGNEmNaQOlKamMraOIzokbKujfqf3kFywvkgY
4vgI2vP7ccqUXWBLy6B+JcDFVcbkWJ/nlUg2bIT/FCWU66Rfm0Kmf8b4MJBnL8l9jBWiC9wOw7o1
+xjjWLgWVcrloGDaiv4y44QonO+aMf5KdcX9k6MBONOV9CaqBkPapAq97AoSEx6dwCZXNDsSf0Om
d5jFYpMjAt1A6CJZphRPa0dHy2NULoBnUCIICusEDy43YSBqiJAGg+3mQyxATewDGyPeXBZ0Rjr4
M76dKCNranKMW0ej3n0ltwU2RP+fV2+Z/TMVsHEaS8Lid3qaAGCHJTgdxFrwO3kyM9nLMIfyXgLV
OM/A+zh4nH7cnQzNgzuMyEK68qws0bBPBqsMow5Nq+Nm3LU9UJmKAQSPGUnwrwcobQOvomL78913
/wfLJnMAmhXjIUUEiHHMM6zAe5poN6+i9PDDj4+ogMQ1UpvkyuKJTUBDFSP9hgUhT6s2fQ7WeCEx
h8FTHEttb2tbvNUyykknbmN6e4s6OsMo1iO/DWU9a2lGSGlB19IG/g5Ot9nuR1+rLTp4Fyq/d0vl
TXj9qCLSxXVCVBjFiH4V4tBGU3rqeSsXBYGy+tjEnwgWGUc2UkBRtcQlMR63+guQdVmg1FGd3k7P
/gL8NYnHGQqBqyaRCzOkjdGgEdBLTF8nXSvUNidsnP4y5FCoNJuvIy8IzrEqoJMmX/JZhiMVfFfk
pxHTcTEunx8UxIV81PwGvfumoSpH8rj34ZVB+bKhEOI4qUW48/ouTd2aVOUgAcrqlE1zAMenPY/T
/X6JYSlDEA00wCbMJUrnKz2199ttntDzVKvSf56nLGYXaf6pt30D8/Rq6nt57YT25noWx4QxdV1R
oPpNnd3CB/udldPmcLNsP8bl43sR9sqjrmiLcFZuBlgpdOQ24HbvLzE+YDPMd9+6xXESaSoQtswM
L/95nFxk2cbmEIA8tOCtqEZy907hzGioQr1Q4QEyXltUveSdRE7GHQt3d/LasgFfTZMTlomCgbJp
oD5hIpoYiFupQ18sxexjx1u+FYeBSZ34b+zvcTx0MXu+x+zp7mBbssrjRrCjL/zdSgnEutjcnjWV
XyDyoFVeRrzR5DPIJ/L9Fm9HBA0lMWKEruR6OK9lbtAL/Bfg/ow/wYOq4oCCCCC0ILkk3U2XGWMf
Mi3d/Q6UCRIuu2w2UVKVmxdeHJK2GfwDHeG1l0/FSvJXq0PNRofFECaERFUgDYwisH67+7nfA8dP
nx4MWpn6k5KBeFCnQnGJ9J+lj4BpNaGSAmpVlDKkwbkhQBAeC4aIAHI1uCb5rWjyfJY7/pJGBF1Y
sLHcDQx18vU7h2DmEzdI5XFUGTmL2LilUD+M+6FYF/ktUTsG6GpZ6pAZ0iyqKjPEUi7XLnT6Yxy2
Mj1R1Kch03/RcNmMMbH/Qo7CGEpq0v6ndbguFpwbb0B6ZG1EgFASZlu0bmdfSNhTGL6LSDCFHVsA
4Anm1H0kVTJ7U/t+Z9/P+wNWb99jroM8PHx+pxplgNeGMNK4wLyWjPx36p3k8r2RCmBH0iAKmYDH
EnGEgbKJm8HboEcsX7Vn2THZHeFgOU/G9bK5KdACUYv1sh0SXUw3ua06Z1KcTzvOF0Zx4kFU3fbV
1oOuZOowZQEeGjdsCDMXv/rKlP96q6+vZZoGVwBYkESNuCYDS96hMQcR5XpBOVHZ/XvbAiS0A2YX
xaX80RZWbtfi0tUFWKHhcPS6jfw7UQCwhVzqMTupc6KpfzCPv2qEJrhserT9U1uN87tW3z+jsbH5
DlT9l7MuvUL0nmRf39Rd48uRx/Y6aHvs2uvq8msdRcFp0IHqV/pS19hSP8iygEer75M9CRHY05XA
nGcWJNlu0195IEQqqqgB3bH6yKBLv6nFb5IXBOkBfIkJmbZMKIyblWkd5GKoGvwnxAHaNWnzDEIh
Ue3JjxrymmcdZE8VCERwFx83zcVeZ8UGgbib+JfPRvRN32NN3yB7PWs9ZKCorYMxrEuz/UBl/bqv
h0e0NMBGyTuuKO43EHBFYuDMwGmuS7VphCj7YHV/4nCYXjnvO2eVbQklLoTM7xUpN06zPzDYQ6KX
I4IkOYjBGD2z7AwmnUfQMq3rpkQtcQUUxs7v9tEX1GBe0B+mJy9iTkFvug9re4gQUFu3oIxb0hsO
DEoOZSUJT+VqgTEG7Aqf/HM74z6eueg89zK/xehjXmP0OkTCwfPTu+e9QUK+YaUKCRgqFdbPe8iA
o/fn/ztMY5y3upWlsNNToiJOVAyka9VoxpCFC0iOl8yR2YKMb9HnkJQn2vS0pPvl5tA8tdomnCaU
SW32cFk+7u2QB8ofaavk5ABY2zQCQNO4+P0mkD7zI5oX3u/uF1yFcp3E4W7ehzl35n3mx0yQptPP
OahpYV1s/7o17W4Vd84h7rrTI/5IJ3uKsIyt8HJWnVY34Js2BJpau2RROAzLPperJRvGaQmGAYZW
uQAsoPULB1kwHuHEdM7ZHln9EIdJjkjZ5+k3J1ZRjCyjXayzSVhvjg1XeWV41TUDqAxOwiS29Tca
ma+PfP2n6qQdC0GtLYi2zpuE4J5iRUxJ5dqEQB2/3GaO8fXfmnTXCEVclXm3MyddjtUUQm+yc+9/
AlV2JiHSfmOfittmUdCcQk657tMo/QYS+/6h2CNeMCsYbxoFCpCGLh1XjCVh1DPsuRRToztXEK3l
nRY+GTAYstgtyozmZ04RQDE5CZZe+HeLMz+lGJ+q2zm1rIiQigEJKLBLG1/+UIHJxfN/IaDas5S0
dNYrSN6lOvw175uvuLBZQ7RLWsW59SN92NzgLIG+Ga+kYyR57r4JO/ZoOv/kjxq8DR0AKz7/4mDY
RHwr38/+8UjvdlMAaPEBPhmwDDVzD09B8knp1cD8JkS/2E83zO2jOpo3hq2Upb0PutSUh9o8GBAs
gi+u1jVQVkSuRDLLPq6/RsgdpyF4zM6s1Fk0BVYfgtm4wK86FCywms2ZnU2JcBKbW3VnYECh3pOY
7CxSX/KxlGbVYjLlvwr5ocyisxbSYK8G0Xw9D8hygcPHjMf/CCR/JuY8dAz4VqLopNA1KgdwtGyQ
zaligNTgmE1lUpyON0MtJ+nSjN91hRrvurAU8E6ypzkpMGDiBS2KBAvlF4mOouFmCrIhCGbWxF2r
SbkgR8ipKdQGzpY4K2aJofXq8M1KtG+ZQ0Y48u+5oIQa3k71gBaIiHcblG8E8gATftE+wcxwEnGd
wGfTQIi6w+s30NaKEMbXUDZ/NtPKhP7WlYPlIirKfXeO0sHC/vdDRqYOxefiXaCXo1gEiQE5OGDG
fv4UnzH8jaN4s3gwXcYVxNczrqYrU9l9dGaLtCuRnPqYV+rcZ7ZbcZDT6I2ItR0jwC/RuOKIsheM
YA057rwky8KXE1xgMITNk6SqYU+qD3BFy/tBB1GTfViaAR2phjrPDQEw7VatG9nDqa3qU8czT3ae
WX+FO2NzsPOyPKGkIBNLvfgjdyZZ3eRCQoURDM/OlEx65fKtPbffFhqHr94bhLPVYd4SHXXdQEY5
j6G71GNqUohWg5ipkrHC92Ctn5L3p3LizJy258d7aDPM6nAf9lnn6fZyJEba5nOEfWdkyEPUGjsH
zDB26ymQLkAAAyNrlvl3nx76SQ2WVdToCziIzyO/QeLzLno0DRzs1WX4Wmbo858B5X9dlRTRmeNB
lYtFc/goXQFF8eVdeom3UXzqWY/qPzCOxQnZb7O5LJx865OTwuOaeBaTl+s3FaKxkMHSt88F8cks
ICFA4ViABcHLdWc+D/yfOW3GdxrrfBFCEXp97j2oaZpFy6ltZ6hMMTpNP6KMzpobqHe5TPed8izc
/WiX0x3xYrETR0LfvbLjteyZEGGrtfRZoabEKTB5MQiNfBlMC67x3ifZzcP+0qtZu3tvH3k7DvtL
WELrIk+WSmQ8oB+wRFnab0yBkvO8F+NSpqGxfTRU6zFqKHStlgKFbytzumrCqRmtBPD7od+m2BTI
QXwaFSaFU7hegtxd1H4qlSsRJT+/d+zCZ7Hb+3g6g3cOVakWu5V6tlB5RvB5JzO4c5Qwjfim1D2y
Kqx9QNW0uO0/1cV2h6UrCXIUnwye8BJBJUXHwyFMHslvWg8YLQqtxxe6CDBhd2A98LNNCweY64/5
I3AQFnhe+FInvRW7pWjUUwYrvwAzynjdsZL48C04bkcMetAtLwCjFx5Eqom8Nod/EkwaKs3wWmFk
OC+s3qF5gfKHFDAZRQ0HwL+kt3Rbqm6H1cDysWokrUh9zcov3it1sCWs+KoPXYstlMSH9MMq0Fo2
JkMVFGYs+xKPYoLh5/a2aahPSSdgbJNxrz8ladzN/KMqwJzynETnqXAH88oEoT7YtnKdMHGjZdEd
0QuF1WMJtSgtbts+Mw0Wn/4KZ78TrKt0MxFvxodU96qHp2MpwLO3O6F8eY+ht4SyIg0AJHVvsB+n
4XWsWT2ETRLwglbsLZpt9SWnPyfY2cIvnnHrIHuAUbs2WokcouUn7mYTb9sFKA+stlP7vu/TcPdQ
8w22xablyiNRrm58bVOygGmW5kvHCATlOVoJ5jknNPa/oU4fgBjFADOmMmof5M8zBC9kQ+UHgfEe
J9W4AeKvnGoMQpb4O82osVae21VuIYFqQmnle23fmX1wIkuXC3eGB71ktX9x+d8HixLNGjFqQ6ii
k5mp55524F6syUD5pLsgM/lzYT3p5SivQng8kTBbHNEh2bMdaJ8W5IUumq5URzF9uXNLMrsj8MX/
R8o8xFPT4YvbZd54SUIK12ffSzsoKVkxWcy9bII15MrDpVWILMdIKb3vw43l0xcULdh7bNmbX8zq
OJKcd+H4h7VvqLlTHNwaoVmt0LoWxuPC9BoSf78i5fIzRwoDRdvqW3D2wPKS8FgtpI+aetFGlEHK
+2tunagYWO4zJRVSefUQVUXoRc2RuWVD0Rd/pP1Ch4jHAXSbh1A5ypD7YID64FB6o7C0FG0KSOJr
sWbQxgb+KyI81++PMjzVHq7LWNav2J8n7RZ8PENehldyZx0EDScr4CFOhNr2fpFn3TvlSPud91IM
lBRsM2oxY9WePhi2fxhWmoxKtm5B3sStLK2KBMzPIDS3MVNSejrJZxyJpb8vo8LPYbhESylXomiT
HP4XA7PDxvV/hIo2CmlVpCV40pyuSyHCvc3ColwKGMTNM3MWUCrNxvp8NtfJQ6vn6Nk7HnXlkMsM
XXy+zsEQWt00v03ZRs6xpg3q5mS7faBFyxRPE5xasDHc+ZXV5cJtNtBZJnDdhiJPZQcQSOnLmD5m
i4KWw2SdlFf2Xlzp/9IZt96mY/NjrXsG9HkUE9tAPxy6tSqURgCJ5g0WWDFNxARFyb4ifIE3nzYe
19SqoCPrEZ6hc24UbREFxg6obShW78MPRfT9kuyJHh/ep11eDExDXvfLOjEmW9s2zMQtN80eX8VZ
EzNklf7hrqhsoD5Cs3vX75ZyXPlGCYtkPr8ICqaL09lW6IoffEAeCSFDKhK0f8aTmB/iEH/mQrsB
ZQVh9W/lL8kYHJoMqoXZt/4PY9M11GbjefU7wUNqIYX8BghrP+CHUziCFQAVGapzkRiQkzWpuCRz
b5ooKool13TeN8brfdzKN0gj0Kg3TZ0d88n6uaFDxm+l4/jNu4r76IkI/I1f9GmIdeiw8Pi8jZ6T
6bYaupniI6PTlzslZI0xu1O6F8VJEwgF8VFRDuLYtv4pANlhY8tO0PoIk8rrkbqPL7mbeUZh3v3k
WeNbfL1E7HWB5LdXwQZq1Dl4/XEB37eCRPoSul5isJrzSUHSA8Db5OjKXikRpUogKWcWyJhQwiMT
ayAbiiAtbZhov5g79RWfNZUZXODRjaXRS/ru77mF8efAlgHL2d87fqez+q7dGPykriDQabev4ykm
OU0jhr7CctiUFaV33BxMcogkHUPAovsDK1IIU0FF/WQzJZ0AlvOcFXDkRD2aqGcPvO2xXl5cdVKl
C9jheumcSt7PzGWgLEN5SVq0oR8hGDZAaBe4wohVbDQoCIP+t5Z31DXjIC8nIA5M8gbKxK2kPlxC
SPTsiM0cmZoKmhZKhcXMZ5o2QrdrsWNi0GXS1JMszQTcrBF91JwDZwK+1hQhR5bUqxLQSOrek4FO
KkgDOafG1IvAzMN/g4m1SNbToFvwpp6XmxSlp9zLXuoO1oXffbjmvvnVygIQqLaZvF1Ct/fLkLsk
kTwvpFJgkRwEsJhALvoAdXvenxMZVPzK1a38wkqNUBGj4BQGgTN8Pxtk+abTyZq1TruJLuYN90k8
b88ibK2AkhdK+rVkdYPUpll9bUPRq0ry+Yr6n5rXo8h2yPZ/njESACricdW9blJhm/jBq4KBVnw3
tPVHMHtxS0jPT/QJxNsEkbzLqZTqcx2XPMJOg6AKBESlrLM7V+dNiG2C5VUd1MbS3Z3ouo1yjeVj
F21YlDpKZgIhSaFlM6j/HlzS0RWtYsjO/iAyEDYd27LLbF7mM0pr6gpUkdoDXY8bPMBJubx/EOwq
hzqXDw5WRU9SJRktUVnjBNVZsmB7burjqSfBudwuUBNM9Nn/EAatQlgR5IZz/EWkATZJ15QdkJIT
lYcQKZkM3HlwYoQJF8pIUUXDz4dvzCNmltZ38zi2h6ZhKp8MJ8Omh/EXWMEA8/+5nBzCXDMrbbK2
imJEHVLuL27tF7Z4Bo+Nv8ZlJZ00/5tNdMzEkaAqc+669NLdbuy061U5V3S3RNImLeY7ljhb02u5
YdKFUVQRXX1k3EfNE6Vg9PXLHVxKsYcV7sDBO26jJSy2yiuCCycbbFK1T3Ssmap8qb8Z3Q7cQyGN
7VGbMl3V0Zi7szfmLJ1zqmYHRBgPPkk8WUyE5aMw/m7ZtasF9kfq/YeibkFHr2IX9PPLHcOTVpPI
q662itYuxmItis/ElBpxmTW7NTOk2xIDYxMpFM4OBnW1I8EVeeaVa1FgD1ZQ1r1XuhFR2D8rbXF9
urvPavyl4buyZona9ceFdZHmV899pDWdwQU2eUybHw6leSMyTOb0MY0LL7eS+8c5F1/8FQtUd6Nz
Ogufbu1nMFi9xH6ud+GyysDRzVgGYXHN3kgcKSBMusmG56N9N+BX7/Q7Gi3WVnP6XBDZcKI2SvPB
zkpXKr8rwF8PRSFfCIhS8a0+9XRP+6WUNmnQf/h5MeBy/zcXW59Pki3/i6rHzGUfFfr9AynYUxU4
zF3BdInEUo8SpRDICFa/6omokPYboOFPTNG4xXY70njuy9Z3X3gx8wWErgjwyY3AFeNI17+Otkrb
4eZiTZzf6o+cZGEXYT188qy1OvovJEKn4msm07KCZxdwCuRewFn1JhJrtVB29Gqb7rtQU9sk9HYK
QK5wFoPqZiudnolCpg9VgvMKfkYhaLh52NyrFSb3+7W9mwNT6B24Sa/J4L0moukSAV8MGzg5/s1B
0T9cE4ykdkgmyO0XIKm5C+CiW5b0+9ixMeYj4YCHVVuWqm+sfjBjR+f2tCFodRr/LM041Jjo1x/V
CRCFUUuQiJ79LJ8jAeVnLjRDzJvTFOiO27RAwImYXm0q1DjtlIzES4ATCGPL4yaiLovWral2GSts
zZTCyjg3O9UNSNyVTTBub3ry7CFznxkGa7FmjVgDCy/EiIwWBfbCPmr4Co8by8k6EoMQIsPv+x8W
A4tRmhiAlzF8hY0heXSusiXRork4DfcwhI+HgiCPxjk8sJ/lQaPfvxkx3MaBOUeOETKRVGidJClg
yChKEuVusivnWXGrB7JOHNIPEYwSvjYpQuz1tD73VZ13Sxmvpe1C7mc+DrJ+7nllwKMKPxFPJBrM
Q86DQC8MeIdY7xycp2noqZdyZXPT67amJo3Vc0jvZcv7u1t/LFnyzh4N/oj1FK2mGS9DYPMbbpMu
GldQuX63JzNoth4YQ5uSuGC7i4fd1GxLi+sbVcNtq8dDDrmQLSNxsual1ge8+YLgpQUqTk1GH6si
Npeqn0cXeYnmtwli6vqSi7mhhARk4ZXlsRVf56wZ84xZ0/jZOggA6KT+AGxsR0IBx7KjEUaQ3zjp
m69hOx7XnX6Hicfx0z36poUR1bbQ61F7mYgiAVaHX5lz9YGoikFxnpKlvJCnJf7n5DmnOcqAVGht
xEDFwRHqHi5iOJZnGjyjMkMSNktdSbol8a3Jf9rFglugnNqVoVOkbb5Pj9OQTwCaVMyQxSNUvFJZ
T4ek+Py05lmeTARSOopRTEFpnx5BSb33k+htrpIZd89h/j0kgX4bxPMitMzNYcyQ2lON6XmKgCZh
j1pJXVK4rUnY53KsvrdQgEgq981/kDcLtsgNfg/0/WiCQnN/o1hShtQfrI+cFP9RFlG6NQGLiehY
eJui3vVVue7ck10wOVmrt+54ORFZt1/n5reQzRuwAKvs4jslkFA1rTL1RKM/se350/Nsb34dCE+t
hM/iXA7I3rvDi7cedOvLBw388VhksgjodzCL7LLLDi0CZU+h4byazgUuUqGL19Ge36NDx6Nv6upM
5Wz3mr8M7gOrOUl/+d3Ue9JmjB+HWd0bD+hMKHx5f61PwGYJ6eXiOCiAR/CLmpqg39URP51S82yu
zDxZThtJR86iiis6rDSObM2A09Qk0XDy5HWvXfYUGOsossU/CUqP3+7Z2X0QbVaVKB1BqfT0yV+r
jb4gLLwUFyGDWM2Oem9lNdwbS/ZOGX3GAhJkNjfOErogutamOo3LurrA3fbuHa45yFqA+Rw0izrp
G9+8j11oakAX15R3Wmf+Fk1bSESWm47weVlheYOIoPRB8Hh9/Y/cTvO698hmTwE9TLZmlToHbsF9
UV3FRbXfM6MCO+6z2opeA54KAZtp8y/cg7hN1SNhJzMqOUWn8RVuWwmz7y9xuk1olfj+giIm7u1H
WeUCHwUgINDDqyGTNEv9UFpW7zzuLLBkg6bXkLUngB/X6iBI+AwxZryD7Qw2lolEQZah70NRzUJp
hIWHjzTF1pCifMg0QaYr+8XUvtS63bQzsbIS09e00iY4IPut5EIAXxCFxkyYgQ+R2Vk5rHyAKsUC
IbZg2VUFuRqmIUsTAh/qgfdSdXBGRASOGH3ZGBz0GnWJw7y9Th1AJWyCSYq071OStEA4FbdYfwSq
MwxbprV6NAOx/DwFSuV7aJewPPTABmKf3pzAzYsTp8OWXk9mrul1LmOJg4zIIkgB1jQTaxXSiaWU
cAGcKPpyLR83SQa3Q5K8biIkvtSR0AqOv0hmBJLhlnZeFjWRZpII450gcIUkiMWlNl8mkZcjEHwN
IJ30KUS4R/L3CTaay1uPkz/g+bz/m7+Vk0E7IhUTsoUlQTWFmSKglZow9blYYTVZfp1ktTlS6SK1
qvyILSXUOXV4kP5OIDkXi0b0ghNh1oXFkllBjAmI4tAvo5+5sAj+V1Q/snF0n6kT1+HQ1kFnqoQt
EJ3hfg9SHvDcCAAQ0P3n1eEe33hZjL9NN02CfyRlrH7QuFkQ2+CuLdPyW7ZjHJwFADUCZ5nRZc7x
DPDiT8+/bg3IdopH6ISptGeCJBgnowFgCIpFaJJuF/ZsBziLmMeLgWikthhLSyK5y935YZZEMsxG
6l35WUSSviYZwALIkEmgJhe67LUVx+H/TjnHws+AcPiuWl1HAKhy4WOhz4m3iVfSUSYgZUfm5+bW
ummv/oL0h2HHfg+GVXzc2fzqKmhba2ScS1D7bhZSTl386fu/OQNSMi3NSQ+7JTKXvRKU6lyRYI0G
djalf11SFbAiZmhzo4s0mpkEKfI2sOWQCZsPOgrorT/8ptIXH1wEIVtxuOAKW4IsOsu7WwGRQW7j
HihijEU0JvyGf0T5KuGsj6JMS9OvfafFaBS2kgOw7/LPcagrAnL8uosaD+scO+oZIK+IntKEfCmW
vDkm5pE/tSAvlauvuhsbWazY99URrleL0UT0h8pzXKA4YJGUT+8q5EbyZnWMPCSC9otROOgpmyGO
UU+Wbl9nUshOAPmCEp2RldmCbiydYe/oT4idpUOQq7p0sUCBBXJAuZO9kLxmAHHVaRrSIvnEPLi5
1nSW1q2INxRBHYa5jxSaCDUSoJLNQ04lRu3rHbdCF1TBsgCjA9CjVSrH77IbrAz+eIoNxTYirSJj
/0qD54ynguS9gzfwLhvYSfe/aj7lgYKikPgIF6SRkmYT0GCSV4B4nEQoZdGVGsj2gMlcbQbvGrE3
tCoYPGXu3DsWfTN+zr/KJQmt4LsZfT4VhTHU/Oz9cdwmkooKGAyET6cu4UNN9hXDVLZ+Akg2gn6r
Aa5KJ0yrF/0vIpQ1rZc1m/ObtOXPVMcRWTCo3nxAUJ/WDe1U4dUuJ+ompMoFnB4cR0ZTuswekjYz
UL+xuPd1A+PIfUKG4DtwRVQ0vLI3NUYIH4/UoTtvBQlMMkR1pMidV5dNlfm0ad+6xcFW/lxCUoC0
i+CU8sWKU15uGOyMQSrEYxfsR8geW9rbcIBr3+7WfkQZsjQ/qVI/ZpHrbjdNViRhBIvLDl8ua1UT
SInVz4wtzw2nhIcuZpbLCV37Es2Xum+AHei0XgXH9DtPJvTtv5hNqQ+3Y/UU8p2F6/YawzmXsuII
qnd1F2Mc2PvTPV8xsu5iR1YdtrAaYeGXmoDRsHZCkc4b/BF4WV6gD5ydDySUgpsbH07Hby9beuld
EPBAK9qffHRT11u9PjvTNUT3YBGRO8HAMYnJv1J4ABCuqICLS02U/5t9VmOrvlOEIAnOM6J2Do9r
61ED5tzuvdy7V/y/m6cWHvYV2pITIZosITM4anZPh4YAmkMsOYIsq2Vu6tTuWWj4UziCCjpyabJg
9vFuRg+SIEYqTfFLpBFSg4L/q2WlNFPJiJKTEzF1jlUFLxyEpmTP5nO7BWerT04LUyCD5bJ7M/PI
azIBIbJpHVR5E4Z+ry7+muMYCPnhMxU1jBC2yXIn057ye2WmrL7ZFxODIdvDdmzzC9C+qj0YUffF
k9es/GwRGFCliY7upEEF6MHl4UHc64NqjvBn/U2GQYe/qRQmyhf+sl8tE9We/L8wVDN05ZreuZ0+
nfLhSvWiLRQ1Lx8z4uCBCZwxLzu05xik49eAOzFQU+eWaEBR0IKkmVu5a9KMvynxufG7zbt68SQd
sNWk6QejlivkPB+lGPfx6zfGgZ39NEJlmYjJdyn10LX6oEW//CM84eSkgVAcABduDPTUW2H9I0AY
agAUE+BSYnq1ZGI8i7SgUsnQ+XX0HmcCjG8iG0P3Cz4Z6B8wb9YwKkUwkA3zr1Nm6C1hFVCKxCcy
ieq7BUZeV1aWc2D4r/H1l/xP2cETM1IZC0WVRdJRJm05ymh8QrGZrQR6/PbmG8eEM2x1WnNtXKEG
eZM2hpykmFyQXZE//DnVqsIXReUO0pB87ELba3UV9FHG3QqloX6UkVqokpeGvMvJCSlogX/HE7Is
en3Nvd7F7n8yU5Oqj7Z8l+qswhfBujCufSUJspcsn7hGvQPgZMs/0FJz8LPnIe0JrjFQZzPwq6cg
7yicM2nz20cdDJ1NmyTQUedVW+uaqwTAP7/X7US8O84rNGED7LvXYzYfK21Mkl5rSUHq3nUtRz92
YgzMAw1wH9mlHEBRI4VwwKm5Z7FWK6cQ5cqRcuR1cVQOKDZbJnTQl9nI9ehtmQK7KKOV3nMAmbN1
I9Ojij6z07/Q2YKx98HxKDS82+4Aer1A9uTXK6OYV2FUpLlpvqpAQ6ePWBmMyRADc0zg4COwD4Fq
g7U8Jr4VFUmGz2o/qzyxlcla0BDVHSNiYlrNliAz96NmQe0fKQAWIFBoRh7pc5UlmUkvZIq8oErp
rlPM1k/p9dBljDXrZb6GSBsiMnrXCOhpmOw7+gPLf7yG32K04GW1kBM0yKJN31USJ0ZsRwRUfi90
rO2dqBCad5MsG9fVf20Ak5CP44MZKpcQ61ZyrHdqaXntBP73gdMqrOgsAtAjkj5QYlUKQ/Qn699c
TShaUl7KTORJEQQfNmGNDdl+PlYwaeAM1V/Zkj7cLmIBamzqkamlfJZACdFSNT/dz1WesJHdFONI
4oB79/uZl4aAucR2YVKTA2nn5ocl5dAVOsoYftrJIY9eH1wTVgSdpMXsLwIx8C94IgnzL9mkf079
g+YIua5infLhMU3e3yi4dp1u1h+Ib8Q/bPbF0u54BhxpwqmkrsaiVI+Ih4ZTLDoKKXE5RLSrqeIj
ZEO4hgJ2vl9MwKzyj2dp5NSncxj96jpqLOUv8ZwiI8ZioN+1hlFeMRlo518qJJl829KDAOHATRLR
ZI/jSgk3GM/lBoPtqli7ZqtR4oF8+869Ikf3vQPaSf0wq+GdEWhYhhLuvJTh9W07CWr01Sl1EHzo
p1q8QCIWWSHclR1LefJzGsanttTUMLBu+ifCzRYas+cUHZtLLFGZ/T1wVRvSRp8JY+YxtBw7edOJ
xPTCEqhQpccpppGwoOWBZoBrTcVpshKRbCZiniuNEAQ0qgL237cPhZjOFXCRyH2llrfqa1hGxDla
FU3MGcCTvdym6jFjuNw+2V/DZo8T12/wpnVVUsZnLuJBVDWFkJlkbKR/mcBCPGSW/kKxNDC2c/q6
z7cKL2LT5BtsjrM+dPQi1MNCRUnajucAChmtDRbNsSAxXa2QbMIOVV0DdGQyfvh1PpECB4cTPKTQ
rDYX0iVIttQiXHwgCnAVCWFg/d1BLAZAice1O8q4SSLMDyrOG7DbC/mN8NiiYGvWxrK7hd9c5Exd
B7Ridf1OPUOIiTqT63oPfflOTuyFwmHDDqeqyXAJpo6i5Y5MO2YC4VqKK6oe3Lo/v/AqaODW5nH+
gp6UUZS/UJXPUaZRAzhUUoJ9HBjpwUd3AiAidGlwHDRofkxFpvWoWpjdNhcwZ7GDoiKVvwrRenTh
tEx+362mbik7kSsa2RjJ+laE+yrDV2k7XF4t7iYMOjaO1bxUhhz78Q4NnsQkHttZmodBcUsW8Sn9
twBFqI1m1HJP2bH+Ul8T0asUnycKAKPHID9Q/0umeDjwUUwPON4nTMP0sKffnmaBt+2Uy6qSGcXp
bU/8jCPfsu5h7QUv6js2n75fXAL7iKVCa2ak9LGi8a1gd9BTASbrTVKNrhR4GIx0Wv/qmGf9wD6F
FpiZuVkcNwur7OmWOsaku4ROfZTCvQWEezj31G+5lZlQtnO/XcrTqH0eYRQlijXEMPkUhoRMB2SP
YkYvE12Vsq8EySTXLng4Y21Uy8ffrbvfWor5WUaQ0JTcA8xM42yViZc+hQBdb39AT5CwdKPiilAk
iIdtZmabukuAJQr9SlrWIsX69Lwv3MDJg/pCj6J8HetQxJD+PmNL1TVKpa4JX+fLhzkbyN8jvFT7
sRy8FgyR3Sib4JYzR5apxdB6CKDOitfHCN2AJFoP/rPw/W3M+tSZl56xwW+4X05ysR6Iw8Z1zNdB
+Os5ObiyoBelWLJjtnFYok5XVBF7Og6IKJMTOBctkPfB3eH2OkIPbrJufLg+sI13x6R5947JxqVe
pQzTNue3RflrmEeUBAg/TdP+MbDr4+4+CNMQnV+d2Pne3j26l8q/eq5zFSeJyrUVTx3liSU2/8F+
5BshdaYqxN0FrO50CW5KE+krp8ftgRrsB4sAwNfIi6TzhWwVfk/5j7U1fvUmCbPf6R19RLotWPxt
XykfQrCctuU6gZo6lgTCKa5A4Vbw0k55/uyDFYpmbspo1gERI8u74y/NG0n6fcNUGh9VCR09yFBz
dlVFGaZni4bu22bbNNFTNvvlS9bcsp+hW9ifcL19ITKCcY9FnKPlQUmIVMDYqaxanfZ7P1PI2pte
zgZDXIslIiyoF0tINHakLkmGRH0NKHuvYGUL3QLG6IysvoGc/XZkZX5z0yIZFAuA8NjiDYYKPPDx
r7AzMTKeJZ6Q7cRUXgru5C4Y2/IpvwlFO1tqn/eft3+WzFH83GASiUbfqPDtoWFbkFgBkbmB+EGY
LscpZQbODtmvu7FW6H426xL7wUu9St1E+ZHK2tvYyD9ntfsutkH+ByBBmucQEyY5zTbKC/X6GMSG
72IIfH3bnm4zlLZ2oW+BIZpa4/GefW2dZHP6+0KFiZWJFc/9R28EMgYEvv+Xvl/TUnYTCjtXkXEO
QrwTvVIVlWN5jCtThM9z4b2bOrQiWM1jl5BVXFAJo/JTEh+cAKT15SAnFz/qMqPctsCJhDOJTsAj
EJmhTG/k79MGygG/lXwoamxXR4xS4RLPNsy9s1pwSofflRneU392HCmfFG+utZ24awvH/CgoLa3K
1wFIfseo4j5vEMR9asIxs4KIdMAqmAb45KIGWGkaR79kycf8bgU+k18OyclbmnWWA70X8G4U/lPI
aoiXceP84bOqYKA4CAGrjw47x3U2AR+BM4AXZleRSkkWbM9C8WSl09NFjqABaYWkRQMMwFb9hL4R
2p6M3yt2gxBTYOQn53pAXhdwSa9GGmXstihAwqK0wRXeahEzmnxcReLm/or+qHzPZuF6HTalAMn9
uIF4WU7D4hn9JfxkbNKFSL7i21aa4q5tUO99dLN7uXKvUWP9FKnwfHjKbxD0hHOIxobMKJDXUNzG
J48sja+Ivn9R9Wpiwh8Z+bwvqF9Kj9TYGba4wdJzGbKSs0MHp114TEroncbhekzr56y/g7orCn7j
7Mg1xJqAyxLyEnXi+m2+b09A9y5CQ2Bk/Dy9Tun6LMApV7Eb3gC8hGAY7CIsSfrPG7xftkqAyFvm
zrNAz5G57mlgblMgDalP8dIDofsWUMuQ28tKtwT39uCH4gq1gDNd0qaG6XMLqprRxKGpsHID41zu
oNaeqq0Fx5GENV6FWDBtV9Jv8EVcj6onF6uYObtdW0+Kb2RkBAXR2NVtmFTnd+e3SLf/WgSTJgmB
67rBj24yqoK0ZG5olKOa4C4QNwGpptCjuecgZTQ3oBQLPH11qIut6l/Wwg67r39wEhEVarBxrDfu
zFv4nd+NHAywHCBe2K++mhgKGKfcJMPRjJeDJo1rKyxkQPQWT4Il8itBk9ZhIXNT+uUj115ntOMd
GgjxOOz8V79x9X0mI9z2E+NBYnCm2CkrmfOu5BU3AqI9ry/ecDN4gLvZOI37mZ/NBpFl8QvQm5m9
gU9KY6wGF3YPap9vhZOZMJsg1NY/B6U0xDswdSR4Pa0C6L6GUe8oKvyzYTlu1y55avFyqM5pSmeu
niHKVIiu7RBjcYk7a7HepOLxzXVbkb5wYrh7ap50RAYWAfJQmopb8ze0mgaouo82BTnG/u9CLfe4
YXBuU6d4WrCuiqFJcIUVcdG390Gbf+kjgBmekZ/mdS8oNOlR6hQPnNrBzaprq35cAncs3GmQN9ET
+YHzATpcFin1LRol4+Xa150XqWHrollPvniugqcPO8m0g1Jm+oNaPgJo44XgbX3jkU4AfyVLZ93W
oxUN/lPs0kxNFabw0f4Rxy7IDudKycFBm45vcDHmaMG4MSg8MmJYE7y7oC/2UOjIjC1SpEwUCjzC
NRVKfhRUgWkp6U3KGg+2fVVDvvqfZ2e9Ne+Gbefla95ujnf5fRAwSHQW+pzsexzSqR2TpryR5iTb
+TPF5rslowzw2nQCE0ue+PcoZRno2BF4KTEcAZiug+2FrQyQLVZm2c1wnAGtUnInJlYYnRsC9mHi
tAFArjollvAw0iCadWNEdGokSKdZ4tqZnoGOVeVGXN7NllhGaanF0y+g5Snb5ZT4QrtP4kBWOFWv
2k7Nr8ZkkRuFe32bai8ccGndmbIwQ2SQJiWOugztlYW0qDM7myJMUGuLzfEaSf4Upy7aEeilPyfZ
K5RMSj3KGo5cGjAPh+knbj82RXAdLEpz3dPUYQSbuy69LvxFB1PMxOWCsu8nyvn+lR5fP/YBrIVM
p/C2fSm4k9k0HxZVt6tEB+SG4P9SZTAmkIOyQSJQmC5df2tdZLEHzz3IxQ3i9+Bt1rIGHtaG3vrA
RhvT1Nesir+96TXU/iAWbBXH2j2BbtngiU7w6zuecx4fYQpCLpcDnarPybjXt++fNne9PrpKstpu
3i5jFNgI5n1Mc0hllVSMvY6rdCDd1I8vGXwaCsnvctZ/AP83epufomgqsD1G88jO1UasVdlzyk8D
p3DWCCMFjx1M1Kyk4Khrq9UCEzrtLZlYDgyGSSfAMTv8j+CAkaTBmmYcO3Q7Jmk4hUC2ODnCrVo7
2rBuzfQjZ4ccCVQptGV+w21c1Fr8amGYXywcCY4AQwvnassZchCBfnX9bRv9PpvZ3mUusIkO9zUx
AxkaRXYnp4HPLvEQdOSM4+OuhG0Wv5Ixzmqff4yZOSDms9LReikRVZ4VV3AdoFpXGvYs+ICdigpD
iy2BR/MluwcCBFO+ycjZeHcwjrcpG8wN1MEDLofXr2/1jOygU+c+OGwFjPlh4MHQHIK7oX2g81T8
kMmQfZptmkeNK/u81G0iuSod7SMPTszoyKVZW73Bt0k1gB9XrmG+8L+7rZdJCeAXDNtPbzz62Cud
T6No8U5pIug5l5AaQVBsUSMljuelZ1AcWhxQjXy3l1NqiokzI1OXrw73qzhZ/X5aYtfVoiq8PERC
v59qmjv/nwtyZuYwOjYc7OFVQRoOU+H1TNEmHj6cH3sM2Q0VD1ru17Yy7xAsk3mK7NGcdSQEF8bL
J/TmwP7hUbLVk/6y9pG4iuhWmdDQ7VrDpTHj5F92OwuLbZaTop+sNcmM6LdkikFGU7/MkUqbn9E2
1ZtFZMOtng26xr8sYSDyiHHe93rHVQy0q/msNn/busT4sWBBqzA+339gX/Qpb84vAVKiZi6BXMUF
EdIVtrUbKNL2+knQ9DbnX56YTl9gZAM9x2Ojwh0goy5uk0H+EwYX77dOp5NyWD6IbiyV4LMljvB9
3nyZFkzyuumlMNK2t+sAvNOz37UQ7ADH7leJP0csnvFfoCy4syOQC7mj9zL8+Ek1qW2+sF1Luce8
vBiTzHjTTZrCbrN0/SdWnZSdX2xvwONCMIRimk7+XtrDpvpfb0H8w+RtEqiBu9pGrdO6rJeWKd4N
NPLqF/SGxFdtKvaFHgRGlf+wGL++BoHaZQzUErUaEcetgCA62isd0VbNzpd23dXUwxEeAmidRD/W
YBfub/noZhPo6CIiQ4+igUSoEHkGXMkcaPMCNHyPqbEZc6MXMo4i667FT8o5lBK1ven/vlJhZ6w3
tDkEr/PrBa7fmHBLF8qA3BwkLnuRxe9ARfbFxrHFyWinrfFLzSLxk+OJgH/7cFhbE8ZIHnNXEnJS
MgMGhSyHMbNzAF/o2qtWT9Rcy1QcTgcq9zolAbvJ4m8iOBt6njMMVuSQh3i+2S1cLHSnyhw5THxe
NmA/XW0jLuiaXOxyFebziL20qWdHpmwLHwjz2GLTZ8TuARJkkGWg6nphc4eFbOx4bumZXaJpGSEw
MmefC9m8EXu4uLLKzwY2MqBq6ASCGwkGS+oIR7xCpU0YTbM6+IV/p1f+b9XZpmfWLqS1PKYFg2JL
m+wI1YGCoz6C7FJFZE6WugXwcg+OIY0wjv2FYCrQHF1067+6TeyOxcaiQwnkkfxZLpC3xy0/AtYS
TDPCOzpx+go9JsctFcrw3PYBGzXD60VWi06A+sKzPRIO90DyLePb9x+LlYXlx+HM31Ivrv8Xi7ZB
/+uDp4LJJrkmNSzpf2+lMgGGilOvqJNAmHyE+cH14in2SIZIYugcOczKz8Q+qnXtA1AKjt7QpFU7
Ya2jUsvWdbE3cSqZHaKV9FnUOlUiz5qgPx8TZg/qZ8UoEZ4ielgrm2O5tWlxRhBaBFes/e1k9GCk
+LGOWxjMTkL+Hl4QLfEJwU6H7ePI6oEA4z4JvoGXmrbH2BycJ7o78RtUcK/a3ieqnu/GR0AuLrLU
szWc/s6+3deJPK2uBgsfPrffzui2Ms/thBGn7BmrpLYaGc+UUHEeGZyjNKOGgyFbzEKvHe1k2/Bn
6RoHQvsCOzc4h24adhoTTTPvSGz8b3v1XpCG9X1UakMW7K7kzIqwwPSK5rnuWdkNPO05kR8NMg5D
D4c2OPkbRA9etKHfXkfZhUIISfJKNzIyLBHZzfRMe6Ay/6c238fdNkU139/zYQWVTcE5vYaJIGQM
ie/rvAs+j0I50A1KFtE4lhZqXltowBZEUYCjCk0MSSqllifHHhrffIm/J0g/sIHWmsRpQT2k4/CS
l2UZ2rxE0dcKNjH7eqj9WU41ePCjCsxIZJ/2UoSss3OWZQjnqFt3sGLKhd3VBWq9Wg6vPfMM4CMI
CetMj/dyU26FaKc76pU2A3sDvu+8LyoDq+t/3VdF5OGu1xVxy+o+G14EyQWhvZ/RDsuj0inm5dR1
05L0oATgK/vFlA89rhy6mvlH3oAN7HcCdDafFkkuoQ5yj+tNoGhcqLAt0F+0BuiuqsV/TQkO6WDn
3AF5Id0PjSJIWOwTWPsxznEZOtHfY2uCgcWRSXwdY/vH3Eci33fJUFfipfKZqdj558/LDs3YlzzI
W6/sKuGK0TeSvn/JvCx7Hbts1HLaBYi6wGIB8epzmmjJBY9rR/8M2ngN5bCmK7mzldfXjcJKpooG
JCIGh9dS3GmKsljBDv683oSour/ZBUM4FZYfewlsSXm8wjtbpYM5+xJ2UCCjDgDLbjQAOeC+Uyc/
ytMCJ1y5q7nW2aNIJaFu1BZZanpfOTPcVuqqLTb1NAYjixVo/sd2EGjqvcpORH9Ig4cCwcQ07e/4
1WXL7moeZKVtUkk8qWGOVi42bA6l0Ci1WPv8xZp22rT7HTyhaCc+YLeX9jdanyqSYMOefSuLKtU1
8WHscJ8/sxsekP2KpzfVRBElmvsX+WzPSlHBoS9OzuMq0l67SpDO9C9YBEcKONeh9SUi49UVW+mb
Zv2j/v0org0YJ1hTtOGcnOA+E2KDlFfxk3QofJI02ktszF5phMxEyr8Da3/7dkIm/PQboZjzTag1
Y7WXMU82T+gHmjMztUbBto72XU/bu0pduIya2B57RH+J04ZhU4MgRfwIpwOtqQWdYP7TzDTDxdNn
lUycOh4nbCJmNBz9H+TTV9eIplU2WBsTb9Jj+FSpoz5LlyCR3KTLVZ0WD/HwCO9tc6hVCaxF37+4
Ld4Mf1mhj+lRYHWoOOHHAQsB1G7E/e6OiP/DSlnyDbj/924UgUVqTKutGB13bFdvkHtkmnmpVxpX
qgM48DPafU3My440u0KkJxDOfMJeo61w4N9vWyFG76D/gceZHDlGFOMenhc7GLET7s+gmbOrmIx5
/ktdm4ggugK7Ot6AmbhjMF5gqEHlui1Ej8QSevivbsADMIBplT2R0rWVIKXbwuXtv8L10CDtk0cZ
zzg5xYhpOk2B3QCET24/3Ea0s4T14n9lo0xyfZqV97y7f8vo3s5doDuc1EP23T/BCapwLgeTLzXY
leVLPmS3Avy/PymYjYkknUz5Lt7T23YY+sSZF8Ec01zow04C9jsBJDFjQeQs2/QtWTrn6d+TbbsU
d9FmFC9r8Puxou0N2yY0lVqP43t8Ng6Wrcy0AEo4WJtdgtcvmYcfuRApn+GRr2RSL8bfqTu4r7yW
Kl0+cwmTSO4IqJtCjh/Wfp3Jvl8/au9YU7l/OqGcnpUf1UNbCNCJrbtZ1t9wqDZStM4YSePEJoEJ
3EMR69m4RUWNHuNL3EGmk9mrgFQJzOcoXvnWUv67oNF9wbFrGsBp+zc+plcWSa/AHo2osjwysfXT
g3y9yt/C/rTXdbo2NlXjL+vKYBQmoD7kfycaMUvtdXskyVV+xW7fnYiExNlScZ88lOcqfQcY40ot
hZF4ifT5j45lGxX/HcYQbJKE0tMER4hiAO5jS2kf9HjATb9qOQ62Uu4uou0SZ907nhsWjjgaf388
sB1wdHKgPbYnqzMGbKzRil2roisOSmAzOGNBQEZOf9hKzlETgmfrpepmMy/jGTT+YAeNhsDMjelo
Rs06TaC4XhcKkEmK57kyhyY0P+pcypKCKD7Lg6I5iBjBn3XovGaJoUGkONSN3Np2Y+GiNI9uXlZk
0L9vcBgmfhm1ErIvXyDwyGuUAM/F7fAoL3EDS3kqM6ezWjDtGV/Q5WnGjcoEC9BQFuB2szVPdBeB
7mThqInW65aGLshcTon5UySfL7N2pKQa19g0e7UuJJhi+0abKTTDLTliXssPnQErL7t+tq/fU2O5
Ht90FzPbrYHNrpV1w3ja616U/BXOzuCayA==
`protect end_protected
