`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gC4Xrgom/AUa2OXRcwvYoiNjl7Gin1Ui3/F5mRITv7AlkkQj9QmwfefWHUapL4azuXwGySQV7Te0
WuXWD/bLoA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KS8VTcEOAbtCP7jvyJaMba+3VO0PU8AuL9kTrUw22tK9kzLzXR0n9L7tyf/26ich6r3lagQxtD0U
CF2UEUm8AYCsyVmt2W8lEqqPe4vYVQCffvnqqINwLOmGm8mTziKHyV+25cpSFiTZrvbg3HLQVDb3
onT1kz8JL2MfrKeZOac=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FKteB6LmPsz1y7byLDSPldAutbxHFstOjTg8CRS/OG1CtN6kmoR89kotIoe7Dco6it4INjU/b2ZV
zhdPDTjXWWqg9XXdlSfFoR/xsJr+bmzi3bmC0ypdmCLsfsDfagWak8A0Rl7o7CKhkVPM6ZttOQm4
2l6My8zSxvao1bnSxCA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l9wEMA5GqBj1Cc43uJVP/nVwYCj7xkzeP+z/IIcdBNPFV0flB1xIrRSFa6cjYih8CYoV+i6ezGN8
m8hLwD8c2tidMv8yWc1Omz9lW9q7OA+hds0X9CGvlNilHAuZA1hfp438EgjdvhyBGd4AKhfvBqSu
0oKSZZfj2u4orzRmLOLvycJ9mVGHZOHDMWMFDoDTB8CL9zM++sA2VuK9SqLMMGozj+pWM1YO7Y/t
h3/sHE033SEYCifGov6HdNQ5ECK32Dz/j8ll8zKdm+khQ3G2r15zkwZalpWR0sfBEztmtVU7TqYN
p3WgcO1W7LAw+rgc6FDXOBn+YAHIKkepKHhJcA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W61T4tXfhcX3Xe17dpQ14PuVGWEFash1FGMp8OSqvjcL+nkMZcBt37t71lLBPmt63Jnq67k85xJb
rKivVi5JsXe11RWX/1KiIeT01hy4gk4O5NKowDtwf9etVstEjsM0EveDo6oJqtfmzR9ngOT3YMvj
LK+9oLmEh8wEtHLLgeGkcXMruOw2iOsT7gATPGJnno9+c/2DbtzyYYWGDqqdLHFrfzOG3lbY/64K
jua3T3EJWrsYzKKLl2X354H6xg/MNECeSu69cbXGCEQnzPx6C4uad533wpwqIILi7p9rdh2Rqvlz
QT5zjeHT3FRR42JwZyNKCBreceBs5DZ89AD8Qw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KaOz1Av4Rh0dOh0/GDOAdeb9zw7Se8p0OyfDuANwRNJwEHSQlRvLVpRUHD67CMNmTe+dLJdIpbv6
DkBktRK1ZetykduGRBahhvqEAgMxIW3TUWojW1FyTKKFdJUmrD1mKIFg6cvtKIPOqSx4Rj9DmOEf
/3trwbiEoukt1zcOXMB4gGW4z8T/tuP+i1APeX+/LrkHvljj+4PMZmwAuh8TNKvup2t+d7CKorHF
L+7wZ816/uvyEYblpttt+8ci/NWsCEmFJ7LEqu0lMdigslUpQJv1j4ga94mRHkRMTBLiKxD2/PO2
C0W29It9IxHHQ9lcnSCFxlrhnQ1OOJudDGqjcw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`protect data_block
MQoQQdmo99hS9pnucsKEhxsH3Y3noiSyu230335hL7G86bks+3WkfkXgNjIExpG4Gfv1bqqEMM1N
3BKg8HudSL2dLUI1pIV2IQ+6KrXbAo+wLTqolwEF1OQiid8EJXjx09z4vbEmHPRieYo8BtgM6iIW
onaH90J3vv/fN3qwShuUicbzp8YWoShqVxSrHJ5n9CUvzHIo6NjU3XD94Wrv02J3u5EwUyhuymNj
kxFNXd1e0NFopvtifiP4UfuyQtz9qUP7aqzfOMeS1eVkk/HPdY8Jr/QWAs0lVzVHKQEivSZSTeje
20K/oI/3AwMW91FyT8ndMvFhlYQOFf4vfzq2UyiyYwpqZxbky2YVVsA47RzAqPWuu0HKAxhQqbJY
e1DhXbezLWqDHY12RstipSLXW7dKcmFIiXOc7Q/hjYspMuAcHi/BTj9PLBf/uKNKJWgrPzCTD9gp
tf/sbt99rtsViHS2llQHK8PiSawCYZus9l4bKjhDpfnF4nfC8P2wakm8Q6UVJ2CEpbj7SjktcIfS
YEn3gIT/WvY1sQBrmNKCpYblsC19QrAoWjicLuIR7AwHrdF1Ag2a6N1iAJFcHtnHOTfIhGFee7ef
mlTnpn/ynpB1R/QfCfMFxLUdnnjeOr/9ZLIwfgFca1/SG8qp6JNZav7IsGfE8J06FP9yZCCr+dOF
Hn9V2LI0oeHnKZbO14L3FZhu8KH/1Q4s4wrGjg3q8GDv8WIGyb3axfCrGyycLSfXR/S+/aTentT1
G7tptOKcw6ungRP+bPmhg3n/WHhhMHTsmcyXvzZFDCDSqynwiIVWQrYrd3zRbBPWMw/y/c9nDrHY
Pw0/M11BB8nNuB1AeEzW0hfMmLcvYpAW/Qg+6wW/drJrrdnBh7dw4pXSTg8AioUe8M7I5WlhcRaK
YJlDepp//n60QulgEx2ib+EsBZNSd6YV1kVR6eFYlqC/U4L+FSOHTwvRvjdHo7p9pl9DXMjhY+Kb
YC6wP7NGuyDUOU/IcpZN5DqKpKjx0l9Tp+6lhrkY78z8WXDKRFXPcZWnQQeQmXaimjZ3Jmklv1XD
6hQ+WYbwOvcrizJpeJheG+HG99FxL0S+8q9PiQexAkeRR5SLZQQ0IXHbqaPYBhfUz70eazwOJsDO
lxEM15BX0VI0yT6JQL/NXEX+fg9jyUuL/u1zuYtGk6TTHmwiLfK68z+HSOl7+bAG3INg7EwXRbq3
JaFY+lF3EZTwq5t1LaFPcAphJ+qhTgLeDpalIbbfo7Z5GeaOEQ9SCNQ3XHdlde+/2LgSQi0vd6sR
mJDKXnzgRZ6t1K2uhRUNMbpHiUfAmLl3x4HKgBhaW9uGg/wrq+Y6p5HRmnkUvE157ZlFCl36w9iv
e6aiHPds4nini98nawNQvvjYFKHhEHPLl7N5GYFhOv5ji5gerWjfECAIKBLTq2PdbbnjDjpCZk4f
48kD2Ty6dwmbw1WAwVVwNHUf7MQcBNqPVFCfnmCTnfr+NpUF35tldQfPZY6s28mOvBkcsJbDOJJC
qinXitSLntTw5xii/xqoIpoX+SG9s629gBpaacK82CLTwxbbnAmfINq3fJ93GqDFz3zNLGlmS9m7
Yy9sDjgpaFJ9W5xai/eHaWFIjtPwBruOBeaBL3vHTHYSR9LTpyHdMRsIKaRSuMHI5Qnxf4bnh9CK
kkAjNrMVOYJ7KS+UWG7vErfo7CgAnDMsI8S8zoRgKKTQpc+JnVPsk2NGkmYUvdrXH26+QwAJHwmJ
YXU5tIlsuqaD5W/o1tWppqsF8MH59JZSC6S1LH8DTjn47g34TetPTHr6E/agTUDgDPEIUdzO/OCz
1CEwKvOAZQ6FDp7p7RlioTozIxB1rPRnHg8u7LGUz+b/tsKLjfivyLYY4unLwR3FeWfIq9lMUWKV
28OMqs4bf7XDwVXeGBLULA6RMK6z0cAZ6M4xYm1w20BDqW29dcGFr8Zk66ioCCriAakzH4lCVnEF
aNVJth/jRDjdhwyprKA5WriBBvOvUW6033pmjvsaEhi0PFtyOrr0mCUU3KNJ2KpzOYbYFpyXITqS
3sDoOVGE/HOJYYE0aWGnKM9Eb3vTLj2LC43m1kZ2PY4FYgV6YiYYt/1JV7VZbaoEQ2kL1/UHCzee
/sBU2gNcLAfawF6eTwBHF4Qmj4aP8c0hVRmx/ZTRQW5a6nLatfsGdvsj9udCZgtnT/Vrn5LNQy2S
tBU50n0FY/42l8sWGpXYrzfkOnpC3jma+7lcedTifVCf7LQolsL79Oc7OBsXuPWxA8Ads2OUTOKv
i794qX93pf8cLx+hPedJ/dvWoI8Ifi6CymkGd2DPDxN5CeV7PUfY5gIgLZNQ96WsyfZt51c5ZiGa
ZxS5IJK+mxRiU0f0gZijaVK9VbLHCyZ6Tx/yQ71o3kcQF7MWY+pIZRj2OlHFLZF0EyUy3fLqyC3A
B0gc3CXv07TPKtoa/5BY6acqvU0BUWeMthIppttOrIudGPF8VmvRk8ngLjI5lvnvmXX6HVkocMRU
8ZsQKVt+Lwz9J/nLLHtutG4YkiIbOwNVpGtuUFtLwyqS01piQ4zgOwU0TJpCpdto1nYreahEZm4z
9e92Lai1hskxA5PnHHZTEbqxXUceJzswdgNrcebwymIojEudAcaeyH3GKwGEE3uNhJcmoJqOleGS
DHcwoOHa3wrkNgRdo873qH79TKfwnnQ1qVqRI600R+SK5IgP3EK/gbieOIAMLN3A3WfuxpIU3yWs
+7oQFbo1grL3Tx3SjhAwkVHFVyj4ciZRycjJRFp1VD2XNyjjk1kGleDLLB1cIiWSCXWbBuv05hqC
/n6LXjIG63TQPETlsP6ohbb+U0IGHlEPKCu1z65pkhTqptzzooeiB+R0pU4XDok+qm2cnEf2+Aki
OWmjXEGJfSY8B3ZIAzj7l3LxvAMOqzDXusQCeL2rVZTI39P2zOI36IUF1Yo/Ajl8t6dPCq8t5kR0
QTRjKkQYqSkwNH324sF+/NBzLiJxz1C0NRP6ePkZsA4acG7nBVk8GTNvnkwTQEUmgE72CDjdw9Hh
6PBswL+sIviXZOMYmL9Y/9oTezXfxuCIGwl4rFKbcNzjOlHwz0Lp6pEdrKiX8wuIpJF63o/ABsgM
2H9nfUQX3dVbRi/FGG2QuNy6qblUHKQt4vLxzJ3ftSd8S+04H+jEjcUaOwOznUVUjRUxmTW+LoF5
jB/HKAqVaS55wS8BJexxnlIEbeXJevJ/5FtRWuVS29IAzyBgs41k0dnqWthdbbxJ12IEWoC6/E7t
c5QIxTmFEMqk1XPGT67Hon5OCYVhYlTR8NrmWeB/1Ytth7+sgET9lGq5Mc+3+Mdpm4VqnSJV9jvz
jggr3zydhEYC4t5+vb2EswftiwTAwzzRCgKsdr8C7rmYRuRrNLuW8ijqReb04GYzPZtSr7z4uMlu
6SrPUr5hAR5HkpLRvKZ8Y6p2c0VxgsnVC/0kOq4N8R9ZoEZ9izBcN5UnQsmdwOcn6Z/OwlyD/0a6
ukBayJFw4is+EY4vlzCIJ3LqmovDvUxZgQgSJvIPzRegsYVUZlIJMntfv4Wov2yCkO8Ekv00Cq2p
0+4Eo7jNOnMFg7xNQkMZaVGdw7fTYsp5ZIM0xOhdTNv1lJdpBHaSOpJMrdtSGiVg9EXXjPNRPIX8
9CsSn0uBPLnwCDxKktITICC2FLSqSUUobcOvVbm5yvZxxGXIbKa7Md9qJlC9Lj2Y10PZZ7+HkZR/
rwjdkxfFaso02iYDkncr6kQKgmMURnJZ+BStB9awUN0eUJr6uQNYXuYP2nw2Sh5neR3UbK7DpDgx
JPUHHYsuh1sK8CmaYutj1tEs6BEUCXECHarD8QN0v2wpDGzsejsS3i0FFTXBnVJ9hGw6Vnki9r2l
51tzyhn1WAOgR2viYa6dMFV2cRnGMpB9M0KYL9qBI/1xPPbY3zl3sqiyd+m2OFtOOlMY+lBENMMP
HeQ3mBxiTsj+/NtawfxdywsjQeg+ldKXTaL+xWM9Wau2DEdvkxXNVdIA0JrXRr8Qvr7CvfiCU3Hn
yyDF6j2Tg6wFsiS5ZsXWw0C7f3UyKj52I65qUM8Pga3uqCMR4X6MO6ikqTiLc3tfwmuyxsuchvZp
aHAVcpuhxGOnW6t5wbG/DVp3LaJm9Y0KZwfFVpniDsnYKJ0LgTxS+nM1qahicWgrEAk1QhknWdKy
aUJpgaGLhwXoOfvSwN6MpZAzczOwwS3E4PH1EfsKmbqkQnnwpOXHziXT/cbpFcMAv+aLC8ZavoaG
8cWoysPg5ev2W5bjqV5IvGgLH/zBV/7EOtRCI6RNYNQG3JMmlHS4qb4ulEHxHbH5DsgHfPRn3b4I
Ae0VgAPUMVh1fQf3YipJqjBEQYkf51H5k9GAKHplh29rcpVMiKsZ8/3QbYoBMYVhq97ZROKiY9MQ
Krk2WGXHOTNY8/o1emJ0v20uzdGs+0+QOytST2n/uFeGpA/LnJlnl+bZrp+SGGXYBF6PPdK70zj+
Ehdr7Yeh01e3dw4lc5kQ6sy/JbkhBww0D6zONeI4ekYyjcpT9e+q4gW98vouqh+w7lqj13PG+NYv
TBEx8OEUPOM7i+iKDANYipLpCibRV8bBt0CduBTUorJrkbUZybsdpXQqAHIeZkmzUoemwXBXGqGk
uuZ6tLieP7Rkq7mfKbS98B8qmvBuBo//nOwW50PtUzJJf0cu3qveQL7LIMfGo7vi1OPXpd2jeAe1
F8VsCHu1GIuCRwWVpqXkrOEzSG4hu+Ui+OtXjUHuqjCjQVCjrw/U53oO6X3UKK5BavJf4MvCUGEx
s+iyIswBuGxhmKz9o8pOO+8SOJ0YSCTPnKAhfOiyuYAt20z/vOdtWYkcLQM3fj8+U/neWSnhHmB1
Tcp1eTb5garoJQZUugCYCldgy4gAub5suN0akqPa8LjJJ0JV4OAaDGIcLE6+SRV79LU1sU/kdGLk
y2sOtZdi3USINde8zILHGn/A9ocHgiZS5+qo0b8a6AkHZ2+z0iTgayzguGP1V7xw1U83WaBdIBdU
jBmATGhF8mCUt80R1/XTg67lE80/oQxJBX4RBbVXjf+PW2fGHhMqFxehsfCtrhOzs5sojPoja3Vn
kHMF/wwaBEAP6VS47TN3hqygAPvXIH8exe83s5bC1waSC21Ys4KeBXGDkHb4Yh4jcpUTeefKI1XF
SMiXAqRctJpDKWIx2mYxtRml1zqq5NMFKo9P/hqNL3at43jIj27QJRmEH9qtCuembMbEmlLENyKG
h33h5e8b7l8TIDjWldGVYx6CKZUkGTI6Ss3cqqf4Fg5O34KwR0shazJ/B79exYT+lc+Sh0DCjtmm
DjiUhpny1srMh2qBlekvbIdwRyLOVgsyk/bcpCPU6HIU0gQZYpDInxz+vQMgyVHJ3AkBm8lsMSx8
u2vJc3SGSVWOZYCW17FeY4CSIILZbzedyT8afcga7p0gP2QCKwAE3kiKfTc0hyJkirGff4Zlh/B/
am3JnBUzYkAQtDO8HBFe+ALyI5jIeEyL4rhjTl6vSlnXHRAzBDulVG8qwN+xD6aNM47nLQUxBkDy
jan2Z27Nvmx76PkplgQXMcKCNttS0kihGIQavLdmR0VO4vLsBL/clvli8pEybqxeEiqKcIlBTZ3h
XEgjUN+rt/edvR9SYDXIPdzhQsj1ZBTxDZlejHOSq86s8hdzOT2nsU8W7NIGNDVnPByM1v9U+gCq
tnZeRhwcexMj2ojBRJTOO17pW7foAvYrXUSxuGlEczxTt6tWxVIzqLXge5rfSoK4MxXOCI9fU/4K
CxeLIpfS6NFx5MLgifd1zXoHiyUaYYpShHnMXIaA8kezW//M8ue/pC5lwPCCFn/wL52BWQbgXaEk
T6HY3i9+kCIqf03plFbwJgC4rxwvp8iVlb+QbfidBGimwUnce11EoZK8hu3g0rqvLuGdSIufu6SX
+jdpN7PRdO0ht0zeQyEtZJ15jr6DIxn+XxLV9BFY62Iy5eOUAtdRbPywNb3JswUV1z1MzMjChl7X
yqQKyLEwcfStkqabpvo06NPIAEupM1WXzgQDjMJwCMZEOjRzyWUw0RC9kVJoTD/OPDYkP/lnZObC
Stb0dDGaqUJokRtkj2HuxY4pGPUvrXTiFgJ7lxnhDyA1jwCYKdYwRxiDNkjxOcuOO8q1x+c7ulvM
AAannsap8pYlqBHspNS7Z4fHemAB0PIm2AkIml8nqMLzU/iShZK4nKsbKqm9rbcgSLEoT6fMIxZo
fLqE4bsiNJAbVParbUXPLhk940sqlS/nnREOUjMVMkpW80bdqebNMJRg92sX0pVQ/PS2wlicUZFH
Sm0VXo84W5xbaNL7Zzm1Uvg5GGRfF4Y8T/edU9uPKOGOnziilQnU92afAlWVmz5QRukgQ9Y5Byl7
gQh22xbS/Bj5OeFBBJ99WUVBOLErXeU65G5eEyNd/1YgoE2ee2hl7ZartSMYbkzWuJ6lTvy8N+a9
NSIonQiHEcg7S24f/sdtYB6Pjz1o/RznGm4ZvDyOWb6hurzZMkrVTdqUwRMSJdF2Vq91j+nSmXIS
QVDiBCyxp8Fh6F/1XVo3ViM195tRD/xNxmP/kOWA9Xw1AB7/ZB45mbxC1WsRgRI4Y//h1enr941B
hD6I0nqM05tTYGg/yfJtaght6jqyfISNu0Sd6/NQzhr92QHI1HnWK02ghLSaCCPAjOAfzbLp6BCY
Cs7L9iqH6CUAQm9qDVwxGWnXMedypVlomJ20EtonQlUwl8abAxkTm4tLyG9fDgx2b4R/JlncEPr/
IqHFdfQbfBtl6EnOGekDLHRIu22kjsOdEBXDxe9Nt5uwWDfDugJhLzij6p8NCPwd9gmGtW3bI4j+
PZ8H5OjzDe+sg7C5zteR09ZZZ/gj5SaBFztKsx0wrsQIDkXwxCImAmvWXIV5JBn7P9ePJUQYx4DP
t/5aTqiLnzZKJCeifbhEAe/nmU3IY3QEvXQYbrOaYUVPVZiYaao7X+x66LuTXb54UkvZ+b0qeyxA
pBOJYICMNxBYI1n9RQmT5nWtqg7I4HUHtrcYBf5cYY9vZj75fyMATflVsf0bn/0sDR9Su3TrnoYz
9S3DDkcQsLFUySkjiN96bat2D5SW1S6NQpJe3SNZZKh6CYJRlpQL7MfncyKHXrmZNJkM9N4/FIjZ
yZXHZqBLA5dk9nEAaPLiW2ed/QovUURuZX77xLDCTNGOQOtAQSQiKhjlxfjkxt3CnH2xlu4moS20
bxagmgNhkKACa/YhyaHyyW5RRlKeRBt7Oa4CxvOW5R8i3QAMeVTdRRpA+eZX3gFCQ2k9nvcEXbdo
bBNshINegoLnaOvVO9puI54FaA1oPxEeifwC/7+Uo8ja1hKOejGQhCqdKjG+zMY74i4IlWzTO+SC
ZDN2RIbWaL9sxxFtenmRgPJLGSHhDTBBTYUXyS+dsOjBakYpBS3PwoH/5SGKsRRp4SqOUlDdVydq
KaOFTGMFc4PazU+QdMfSQc/NzrKFX4+lYs/NMLSHfxUGYgVnTJm2Hgg560CP7me3iNBsaXORi1H+
s2Mx5HvOVbIsq8wSNslZ0iESA+HTGsZqoz7suHjiYQj7jLPqBUFV4PQOpeTXTCGJNaR2JA7qG47T
yXICMCdFalciciUeDEcNTi2E3SZ/8IfDtXOg574AuaiSEUKCNaR7XkyfL4CVa7RDHkoNVTck5dnb
zqKDv4FOVpDP6yPmG/0OoPbIyAkq/8WvZw4PRauVrd1C5mKSkmXyh+E5sM1yrBktAkr5ImyHQ2Tj
yaeOGklJj6l74Z+/4rZ+PPFVu42VtskFofzCrQs6aDe19bvLC5XIgCQE9uHwmWlH9hbxF/yy3pc+
2nXPWBTB7YuLumtJjk8b/t/4dHPKe3ch+ZrHCsEKKEVRAgGVA9BYE8r6KOz13ZecED5oozF4eiOZ
CyVO5NmwXNDXCD+xFtj69OmzbVd1kk8KaScDDu/pY9YWTKaiVdWNcG+cjShq5HU1weHWDAdHOuJF
SugjYsOwDP1rdm4LRtVnfSSXkjsXPeLlCSQll9kdPqb5KuW863kifaQd43Me5lnaOyXmggQrD9fu
2OhbM05UgKlSIuDlVQbrfQx7wVoPd6zw6dklTSRZ5YPilYNcX2MFDyTdrD5vHX0EdXXO6+ndUpdz
+wzNelwI2tLVUyzQvlHnGo6me9frJPuIj10sneN8zGtBymeW0RJJ8EBmb6B8tHHp1/7lEhwOvAEu
PFGi/9c3SlzIg5kGXWkrhjFKv1CZha0aecoZNuUoQ+DAZtgaTHz0S1gOWHG8srhdpCARswDzNi7w
kzc08PWxvfjpSd8+/QWzN2LQGRwTQKgyTZKvFvatQxNTgrikk2xVYe34pHQbo7r53Dyxgib073M0
BIbakfae+494V0BcoLW3/OcdECgeRX+S5VmZAvvuPscJIexUJ7MhdvtXIr9OPTwGX97dGpcLyxJB
GW22CLhmdkVKoL+wqmSNUYTfFkfqxUcyHuOQIbLoZqXUQ8Kq+oznFPkhPk/9kbzU9eTmfkkFfdMt
2Iv+QenplJzQshUpUQ09UvuBp31VPtSTRXFRArpZZgT+WvSqFbxQATGlCO+tVhz3qc2OFiq5zZmK
wf1tCMDe655p16eg/e3vFP5Eu1seg90+lq2f27kwBbvM6g8j0kYWzHomravT5GeJ+phgSWzkBWE4
AOFseeNTvW+srbGws4iElGHRERC6ZHqIC8jDV2ekP4AnmY5YGqncaiYpY+lJtf9aivk58RxTCBAz
5qKIxOvxZ138pLXtlMV6Z+hi0HLq05+Nm+VaL2/7uI533K1hf22LA7FUFtnTipR97rWBL99FePah
5LC+PyH0zcWoaA8xQ0qtDxAHHxyth8dqgAAIKEoIJ664e/DRB59xGUWRPWaZMEGHaLV+UNfHHm5n
fPX91c7kmTpgZwzzUC/XOhQNMuLHr5NzpsDYIrq9l3wKV/BnRyW8SZBywgzaMePiBrJtgWE39/e0
F5Z04CIK+ue2CINZEoVSLIshoLDMhJq3Xu7Zvg3X956+Iw1Ujmt7iGyd/Q28p1V8CCEqhck2lj69
Lpsa0yTEx/bPcW+PQYvtSfrwYCb83bqRs5l1OpKzhKP3dQvzh7ODQqHGZmDZt3for8DJzWUc/coG
Zxjtu61GqQYWrNiPPJKOsbiF0qqckOOktZ8aCINi5hGgIHy21so+F/yju+YPKFPRrhd0rMXtHDqa
z21ZZrw0Fp1t68DLsZdE4Sb4HfUpUZ8maTXZfshRYCB6rhjJwdGYBVKcs0SczdZ1U/rujBSis3o+
OobUzxW/z6aIFsdLxw2czYZek0m6uTSPD3993EU6vdoIrKuAEcwmNrnUpqlAZMJOK70h3FThmYi0
7ec2nuopsW3Odkc2VylyCOv7WlvDAxUBrOR8GJNINf4JHIxJTC9EGxfSSo5zyrEoRDExvbD4lniw
4KOFCH4SXDyULir4cs2EeSX5NUBJlKxxiA0xC7o5sVbv3KbT2xwbFc6c/DApTEPpSbSEZCqCbuo4
gVEWWp4LLJVbDjltrlyhWleiVtt4exyT9Z+R6hfJR0rVsy24wybxVALnnNm5KcBtauXhugbLEwSd
uTlycj/h6aqBIomxAqsLEAmO60tYxHveb45N0hYPLLh17JQk6lqeYwfHYuzRkkXawmcNyqicgU2n
dR5SB5dhf+wn72GiJaMnJ9a0EoMkvKfzRZr2RkopCgIEqmNH/5Pbn3E47dgPuapE+REdh/smDdNQ
D9xdDtN4fVjnvWu20+85jSp64G0orqACilA7lqpFpEEOFXI2UMYjXWLTyHLFKFBpdCkGiqpQ21sG
226OHSraGhiosJy5JyzjsqWeOfl/dSkdoKKWvTQhnHIZ95DPtboQIrHbxFu1qwQ5XAAEGhIrpJTZ
EM/Pbe5Xz5jBZuFUQO7nWGVicwAnVlWjzdLmzQ/fw6Zxwp2or6dqegkkPlEpjEuoMnKbNTMReNrc
Sqo8XzjS1BtWUgVKvGZb9POvTLGnwvlmpFogO2AA48JvP3/+HbaKuk8K+MXUEadT7cazBLvhObgq
9u1CBw39kvptTaaYluGgqTIHbf2h49blcP56ZjOyaLhoqePuZX8v0+YPIcujzNlf6ixI5z4oHgse
Pfq5XrQYr87zfGU6OQWcNKJDksqP3F45za9Mvsn5YmJU87R7hDJKzDpzN9l6T/0ic6DnD5n58z15
PVwD6RAriVILRwodfnyE15j8U3WQudIWfL3ocS6Pwgtt2kgqRlTLSgCjh78aEHwEwyjZ/nmxB4Gq
C9DaYZbcWoYagEfVRKnJnZWQEnFMfr2ndip9WABaXL6r16EGqCCzZxWhwqlYV7Mx3urR84xnMF3q
5PQknxyYO39mULap8XaLOPAdaFWJDOyIZBF/sIoEk/MdklrbqD+JBGM8TaIfhIkKfWW3m2MgQ3DT
b7FZkITJMA/QBovz+CqfXp+3tphKz5VD305TREHqFOK/syRb+IX6+X/YPvl/9C24iG5WxUFthFFo
ykQMsNI9eDR69CUcfhTD2QiF1C35PknV1Rxi7wLZpcTalG2mq87T+41afbWiF9qnSZ6Jm5UdUDLN
dYoWEStI73kgOkAo9bYZs5WXDJBFeFgomggRtnPneUtws4VYmVpwOlakBF0s9thm2fsxJzqW4trZ
eGelZgErUD/+nfJXwddQ9xoxjQtE3vUoQWRxbqr74ix56PUkHakhsjJSk+yztTBOVfWQHZgh2yiI
wuofiezcYCNM8aH9oDs2d6LeZM74iFoLw+6DeDnRUSAlbDD5R3oH3TJm6UoahhkOv2CFdXcWXAbL
L7jZdi+EREnjkaAxeM2fjAjsqJXigwgIb8QPI6rXY/uLhvfVUReSEacqS/u+BbtLr4FP6NDwI9rA
epEEVk4GySmhW6VmYbF7CasdnffxGTAixMlpQ7BGGwZrUH4dDw3VSfKcFJYX6zFYaZ1OaWF6gXQq
vDycGGiG/qtACtD5c65aYuNNI7WbCGay/b5xBDW8F+KQimMEW8XVkYjGKPFonkNtdbPzqi8L7jqw
tVuZnwrPgd/qJIiCXcMmwbhCUYH8LL/PSI9u1RKuELfYIEMSTikp5tiTtzl95uxKkwoN3drKjJ3M
OKlXjCY2Pkl/S4n7PNnSCvzz16iR1irSDSoUfn2dWCD4nWC+fzSncedNSmoooS5hKCNzNApyCyZE
xbxxzyo2gwHwM2Mn0Hqe7908PmLZCxbmkqzbQgHmmXSAhrVcaSVsHpdHI3iqNgc+M4DHUJ1CKR7b
gf1R0IPGNrpfELSE7f1DgMgwYDctCDcy1WUDtVF7g0nYXmvRFK+fM1F6fJg3gV57HdnYsP+M2zRZ
FM5Spfwq2ul0l7HMlae2oC/SRu0GJIXTnzg5RKCQn+dJQMjdtXVKq5L8mEnN/Jwm07ODXSs0vfhz
r5tMB14ipBMYaWGar+d8Dbp3YK9CY8HPNTMjDxCZVvrSJsJWja0pLGmNipzFIDNb6xyAVuUrZ5qQ
Z8ymEejEZtw+HA4iHrCUUphP/s9dOvdqo0sbMfxrz8FcsI3MLyiPn7JoSfKoe+KxEQJtqQz9s5k4
uj/jAALm8mFsDMOrSXbAGVstjXyxtQPvSVjNj74akPKZkDaxMmxhBeWjbv2Fp94VcjV59Slw9M1O
raStXbKsWDhRLx4hw5itusmfsdgaz6R3BhWfYiOhdFnglURcruyyY4rIVLOPCxfFpotw3N7WXLTd
BGITp6yoNBl7gP+t6c1Z5R+I0PjbevIDbb+c4/syhAO7Ks2FGto2Yo2rjzpuOXv/yDmZP5b4e9SS
5RACUlu+pU4LLE19xi0q3IcfgjttyH7DQdqJzRyw/4pToFXDY/uyr2FqipKwvvfVvtWw4RBS3xQw
madDouM8F+Zj0rxz1MeV+Vj4tcdy7lynczI2cOkUdFQdD1vB/RRC3AK+aCpym3XGdJcN2ZXSWj+M
WNJ1V8ebDtWOmY5E6m/FnO0pq/xpcnOLCrbrJBg42InnapQZRPgrfOLzevh1wY/0APPUlct/pvhT
FK5uMTfQdWhN/TfMJutjq/s9X+5zxk2JdWS+xfOUl4DJ7uwqx57CPuaBg1DGoKMBuH+ezT79mScW
tewCdEeCwYt/7basrArnqLE1u4hz3aKp4+ywd6j889SFLUbDYZxsPmAVmKIsWELt43M1Kry6GCZi
F5x893d9ix1/5IsKA6bb5EoyVH8w2XtE6FQnUvCiQoFlxcqQ2uFBbvNr+DeLOwuDBSu4dYoanOUl
3z7M6MHO+GMByGOThPhFdeDlDhGcPcLVqeqcITxxTtQoSr5UJfrePv9f0EZDlAv5NQkNfC/4yS8O
JZtgco8n/dHX4cDTPyfmYIeHyXlUUAbOeaaZ+pwxQzeGo36Fip+tdPnNHVd/ul5PLBseF4FBpNwA
Us2Ha/J8sslV4oURd8woIXchvPPwTSOe/OXeQhpOOn2pVS88vQF/Y5WRKSDK6HGnwq3gcNqYnVRN
d07GfFOP2Wr7wtpyoHwK1AvD9Obi9ywkCuNjiVwgI1bY/jySdEgpw3EN4WKomCI0Mi0kb20EHfI+
SSotBZ/4je0DumwWoEjPJS7wTZfMnF7LYrkyQNw9bQOHxcM73yNcmbEwBgk8B344DGwgzF3cmcFW
w48a98bqZIF3ijASgwFvHvm0gkJpHI3ezrj+mTg7Yg1+7N7f6VipTxJ2qcxydyoQi0NAYrUxjDdT
UfPPhvBE8kR/5jp2FSuvqO/GPpfdULRx8x2z9OU/DxuOLbM0wkytwazxXezww/rvBw41cOHHmm8Z
dB3LoEuS8mmcXZ2PSjbRZNxUy0c+BBp02dWSc6TxaVmuVpT4mddUhVbgd3Ks91xKOZl9FPSuOYmK
jtm2pJpRB6gl1n32U3M2TaJaze9ldax3lAqSa9wjfHFvF/we7HGlawQZ49UUIBl1GXd0+8wm0z2U
xZ9IrwXxLF0IHChNDelqpmqY7CWYk35FaSBDnTFSy9qEiFSKF0YTUlJNeGBfrw9BNQmlfb5sxMRX
CnUA60pVgf2l4kNGUjdrLFV506OojSLYoiYcydl5y6utD+nTqEdPQZiZHS+naIEp/droV2bIARwu
DMx+mEwIHEKHZoC1LV0sarcdqiEFrhTdKkMR2you+zCOA1MlP/XdH4WrvJv+2q6nsvw0G8fUUUIB
pA3u2kGlMNb8RXQVXkok7+l4vzQrG5rgGJltZv1lW+V6Kear1NrElbmYt8IKNkIKCfLJqt3Zbu/t
7xxFApqYoMc2sDQj+itc9APKh8lckYB54zdaUm47sqTBdVcAzqEnRaqbYJrE66aYWnGW74KCgfp9
eQto/um/ioqTqQ883a4W5MyIUsvfdwM2snh6wIDCo1MbLka3t9fTsbKhuJBNPRA+W6nIuedrOp8y
cdzpCSIsuW4Bsx7vvzJB3st8I8oQpXUl9p2emb1zDv9Bpmeh2eYGNbOQmDH0Rb5j1rA6rmqOugWm
E0iwjLAbClaan9qpg5upeR0+dddEFTY30ui8cfoahx8DFUOR9aDiLBdN4NUJxsSIm829Ojmr6DBB
v01jqbyqm7NCxlyhrRCVxRbgLATqYiHgsgSj441Bmr4dZ93hyTV/GkqJVuVZxaGkk9deMOE5i6fU
6ATk5O78DufiM42p24s/qf7LJ6WyXE+WCUXQQSA2lYQvrl5mMmykucr23ymwwSHy5NWJCLEe4VJZ
gubNfezHp6wVw4QSwFDlBZ0VRxzHWINXCcMglNBZcqdf3a47I2yWeMAFqaCWAHDi2ITKFI2N8hEY
3mcXN4TlAEtjO8KpWB/885Q9iGnA/kukd+ca3cO1m73DFrAq7sr0BcZwMen/a1f+bDZx2PnerYvQ
nDrZZz581V+EGrrx2hoHnPHdcBELVNDJUvLIkaXawFVdJOIRbfHXnfJVK8f+0rTlMV3XOKLMVx+V
BGGxGgy8Ruqhyg8kyTDlFDfOYI0KSnF7B9hfpFC6llOPXKmowWByczSQMgbk2zakDnpo1YqPQJF6
DrXrDJFAyRV89V/D1YT133EjgTCi37GVmxdwnhMQIjlNtJBrNlF5XTrNPGJ3koWSyNQW3Y8A9xZn
MeDme5e71ePaG3oHv0T03LRAU/f0FkWidIK1JTm5qdxE5G/RvrrfjGHaz+rFNymNE0730WJJ7oyz
FI5NuLF/R2IKmabUsKaGyhP8WZoEjA1pgpksPXml+yfk1KU1NxeFJytackU+cTe5Nrdy+8eGfPch
JjJTc5fUVCXiKwcZcoXMmvT/PDvVcart3TJnRpAS6kzo/VjO214P7oqhtuhJPvhk9+Bwp7PyksHB
VNT1hjWVKHyk3kKWEeuGm/Ipz0VkbF8dagpdJIrcfyz9kfDbOpDZDD2uEDwQca4lC7TOsgt/zyvi
ls2u4qKwiOmlxaugaZthPEMmK5es4qawnU3EcPCVUzLAlSTCdtIQunCS00WOP778TvfsvjD5zXKQ
5VC+v9E6ET0C1qjMTDkhYBpgvwNEI8MYne9ABc8octPWGD6Tyso+8VzGLMfQux628jAbCxar3ELf
nLJ29dLhWBVLJjt6smcKE3SvwGLHyxGrq52dYIwpjEpYi/KSTZ+d/a6NxpYPXFAPAihP2180mN/Z
2ecW/++EcKsTIQqX+BB9uVcUZlLj8vYjla4XHykoOL3R8WKxUN2qr6D7yjkFveskzRX4YoXi5owN
ZCetC9mWrX4zt7hHtQ1DEW0ocZW9xj+Q97kf2In1hxOrWmF6oy9Y8y+tMBRj30J7ifvQvU7QYHSM
b8bdGwW9pU1hg6Cp990QD+6XIAJ/VhcCQM0qjBCLe8x91dMVMGsjBvjrcy+QgL6PEn5pUOlavaDm
0q9J2rEtKGw+kBebGcSXYLfr4CWfF6vI8ABmXljqWp36biYpVZUQ1JGsnKCuFKisiD7Vlv7IkCGY
L4iLoi2P0ZyPWFayFll5ZGXnAHiuoFqSwiVMe1o/0SjBM0m21Gdwwuzrx0KcI47Q6uOOcrieDfwS
0G/fL+NVcqbtDEQCHDjiq7LwRvRdJ9teP1IiwnwyfLnZUzAOYPablDIric9m0vpfbAo3t3bXZ0zZ
0XI5TYJS6WwzM8IvKhLrIDTRCsBWllt6YYzf5D6LOxqfzA1/88J+xo73Y7vGEBcnqFH0OyQbEUDT
/0KpdZi7eZJXp0s551UbQa4RmNOrtopffSQuZdN2RxyM1SbQyxUonKDPwl+NxG8XDG6i+PIFJsIN
vL6UnZ4bVV670LeEr8vzuyFFqNjOqoSF93qxLqqwA/l12PCK8iBToA4Z/oS8/3J7zk2iditkjbDf
gpCvN5MYxJUJHU0vOeth6j0zmp46xPpjE0VO1DcYj4qPOB75JHPEEInoP0NLPCc47n00M0uzhpMt
ZZPYaxQ0EDuv+Raa6+J8b8Og1gfC5d73l24m2OucpSjjWj2wIp6mUc4EQE6FNso05+Syjk9iimyN
OxgiN4sJ9j93BiJDk5IyyY/knMoubIM9xnZXYKkt4Oj7oscWAQ9H2oHHT2D0puI4nu5QNjVVWrma
JTYt6clRXzQswKzSuSW9uzQD18c74lykw89GTtyVB+yfrNinOeW34mvwS5ORk2f7ExQGU2fGp5Dd
PUXvYdnbh6FFevsjVng1EOPy1THGWwLoqSirtsNIqvVzIx/MOX4/V6Civt3vMP/su2bDXd6vFF2d
LfHH7vUOrnHQjFKhBe7uPfyKBI7rzqZkArWW4jWK1A27dpLkw8MW0hZvwxL7moNYeXAxDOk76d7+
SQ2XVS0XZ9FcU7+jiKNWFo4B1YTS5TWhTmhMfbFkMlrojEAUZwdcP6+K7Q4baQTnPptJm8SA18L4
FozbYHKrC/2A42vGXp6HQaExhcFCxhOrl0S2VwwhQ98h0y46rGNgvz01fUIu1Dwm+jH0U/SFk8RM
jiFASNeblAE9F8i4rVBsP0E73lO1jue1cK3lZ703hC7/WZ51yFKYpPEbdEMFrRiLaOskWQCin+Z+
masN3FkPrOo9w8rPzWVGe9T4M7dWTSuAxo0NWZzFcBUe1PC6OvzX8ATQc8vA0dSAmLWdvGixeODK
8ov40Pxm2quIb9CIE020pVq0yk+wLUxU/s8jpFxts55yXtxDrqfBdMHyQTh54XWcWTt0Re7gNWHB
vTodYy60376PJYrzsdXKqXjFxeGEHc2JUyDC05XAIi5o25jq4zKt0js3Y6ee7NSPsZ4zaH2EDFMh
r+mIAhdj1zR+5SzEEhikPyh11KYn5cpfW0aM7crmciKKX85+8yDxP/NO+X+CGI2RIUYY7QeM1ARW
IWxlcnEKkruGqmLZ9n7Y1Ze7qkQmO7dhZd+hPIT+xtSR+EMsYjKHqfdTaKxnf9X4Y4acl2iYQuc2
EDm5opHUKYPdr3v8KfMGXNuGZa2CvSv2nh1AttjWPJz7FGfh/XaQQ1H6y09dCOlnA/uXHFS+9Wk3
VLDxKp0pf9duXdHoVMyikHM0SsRiwVlDpcPQ4Jw5xHEA5rl+WujrJy6i8i7lR+jcpkAMnNgvIbmI
OknzTaRZk3uQcw0szQsMwbi1NIfp0Rs0Eqz7kR5lpdVPCuW5xJJhR7GVgjIFE8sNEUxWy7p3ZjXA
WH5oFXkybt3atm1mP9YxIFId7f3tFNpyHLuohKVkAa6DuGCIU79c5FOsazwRpMGxrFTnFiPGn5WE
ih42w8aLVg4ebfnphVywy1VfSaWN00rrEakSksXOX3nsF5Ddg64z+xMaGkdqH64CZy8AJt70ACvx
7qpHg9dbusTXULtyjwg3x/6y+o1bO7IWc0/bCzLe7TTrAyPd/J2QrFCdTDJLPg8u4P+ku/nXzYJ3
p28yZwVLOtGwMf1GFSRJ4Fo+ebT8qsT5po12uyaID7+/C2Ja+JhFN4ovy7wMoIlJyhkkFMw/evJm
YPVvUjAJRcJVFkQijqzEA/Rbtme0hVnn+4UqfNlCbxA+2LBNQomm4nedny53MB6sbTkf36E6b62T
pZpWHmZzo9XK33PMn+VHHxD6KNBmaVZizBZJkW1M7sL5Zut0n3OUzjfJNAV8Ao6YLeMbKRETpGnU
jP2zNwH+mb+D83m3USHOOoZXd6NuMNpXuiH+3Nt/H3TiW/tQ7HodFbMmuEeVwFMUzgHArH+TAWls
JP7fOrPhfL+G/iPPl/05E8vknA+m5FCfObVZaJJ5gA9gngpUJvnvj9HDPQyDbNHm42omJlbwqobM
YmWoGie2QOGhCHcjn958TLpyQ7U2On/7O6nU6WOGzE+8OAjFAJQjTemtaEI5apEBZlLVnJrp9ccH
DFvuCVCcXRX4EcWqdAWsxXvfCoLsz+phFONJCVQYauZzQs3QadQV/NJ2KpnpnxZJGVkCiJD3u2lg
4Nj30SYAGbM4VinMA+y0f5N9ljz8q8xtZK991juuGqEvK7c4o9rtMMefReFkWPXYXpRsBYf7YP+t
HeMir/muhXHY6kgjgY4cSCQXbYDiaBMNkZ/o9VvqhYnOTrWlbOy8f2AhpcyLqNQklpGNZUyhINKt
U/YuVlRfx0f7NHuq4tQs+ma0+jJD5pwIXhd1GggcOhYEokUluVGkkPHPMwj+zrKycdVBv50tqLde
PsjJvMkP39k/fgMIilArsUgG5Zhe4hm/roAUmuhWzomHcpkdqIL5fPlZWvsQKSIWNNQFIySHEtbV
WkhzRsqfNrsSay8pkHzLSq9kUpYVrWM6HL5834ajFgMBgsv9QA0LfW5HFU5ojvHVYVtb6xl+o2Xe
BxpYkbazGZTIuvL0K8XX4e84SXyEIXO6j4XpuswZ5jxs9avLwHVdayzbY2oNF+WifW+Zw3uIgmLN
hotja5H+MEeW7PTB+7ALORt4jFhpFnNrRJlnFKfWe8WsScgsQKJBr+J6IvW31oyISdzeAaicABAT
PbAMzJqXMYHqPM3pLktynfpPXIDtsUHTS3Px+C8byEgzq8Thb26lOqdoLxHO+DnniZsmU+T/RxMO
tTRkqoqwbz2v2vhGgTyxnfyOch3sk7vnjFL5+eFcyj/IDEK79yAxRy6OhkpRPMHfqg9NIX+nW5XI
T7U1/zhKph/jKJabYlocFiMTnU77IHHecoabsxoLD5lFEa5M1wRYdgMgvpljitpt3zfup7zYZReE
UnUs/Qtj+3+nTuYWAzDEWm/YxgP+zOLIqeVFCun6UnyEtvwKQtc7Nr/5RucxkaUYp43gVYwPjd9B
CWWfUYu5FYk55xBFrdZVaJfUaSQmhGJsCpoIjS3nX2zPTfVdrEsZ5LlT3Oj43SfvYNopax6dSx2w
0A3HoFMwywtfiOmZcMMj6fVe8hHDXLG9nPGd/DBJCdsEhrlgWtAm17PuWXgFSDmNuSVgC5XpUb9W
73nCGT5lu3FrtE8RcxZBPGWBWR03JfxZNZQJZ8AzMIWcYYnjhFR7x3TwzFAF40Y5WeuAH+T+JTIu
kKaYRVYMsf/gSb38fpowwZOpngjphxeUy/5HSRrgFZcMF9X0Dgt4i4oJzOggvwwC1P445XImIm5D
uG15bcVKte1JC3N0H7g3glLSD+677vQsjOT6dr2Lw3KqGsrsmuCCP5q+VhfiaCmNtjHbOt/d8pXa
N/CV8+V2tYtzVeRKKE6AqIkwzkQwklXNjdvo854U5AVqwmwuZK5vAU+tJJru5e/KVEqqlTmzCB+q
nZFC34XB2sR9KpXzaLt/Z8XPimAzPq0Z5wpWSuHTRzXp2hmYU//DSxQ8T1uUeRUhJQkU2GzbMUvE
3muT6g6yOIXlFrDZPb07jcoMMeiiuMuNeXfkpPQQ7wq392nLM9jjIsTMjzVf1hymDz3Y/jb7QFX8
B6p7qMUm8m2JFJdhpbZguVlejkrzF+zP/lqbimEQ9jylZTchbVqBpQGtGihvnW+ScxqVNSjuIMdh
WPStZ0LftS4eYY9dBYU8QvvREBbf52/mRlqefOPwrpHQOeLxnBbhDHBcUH3QEc2EM0cIX/Xl8rrt
dEDpZoGxNQtrMtQ0P4Tx4Rz/gXyc8f8pN8XFbK3s8NBTGLW7mni+11xma+yLQ94KIVVkI7haCs4y
B8VARwMFuCOJUKSLQBHio1gynbb3LfSxYCgcO/BZVfoWCTbMlQWIuryCnC5iqda22B65memwymTJ
5mo5iJNfCH4Rv4laV/GYqOPX4NFnvLsTj1si8ic/nDIZXMNXzweEuZ2ZNuP02ZoNM7n/Njy4wB3c
iOsQZUlnk6bLUAOEjIDq1Z3739MxMS2zOyKr7ZqvGNNSexDdh4JTKYMvmfzJlPTanwlYfxKGLD8E
3+/TxXe++927Ah/N6FL/e+avuYNlh1fIlTneVnO0A5owLeJ2kqSd/cGiEM63hVRh7zt4EvOebpot
iuV0MnrN79GqgNH76ijzy9732/T2ZOXlZfdykqAN5gVHjGfjVM3sOnhtaoyHoCr++UI1iv0Epq30
oLd9C/PdgnaGTfa0Pm1YXfZs0KU5iEQXjQ4Psp+aXsEzhuHY98XdyzadEeL7hcbSEEHWyvUdYe6V
3jXUDR/zsUAmFn8PY9WkvGesrhCfhsqGuVm77R2oHnQ7Tp6Inei3k1BbE0kE7esoJ3cF9TWqlQN2
m8p295MK/yc49Fo4w7z9CPC/a1KnFljdlCWiuDSqBfngxlWWctO9Jrqgp3tcFGfE8F7+c8dU+mRE
wLqxy4HwS9HNc0ruk20W3/3/nCk/fcpGL0aG5CIzvZ2ZHqW5YZ4BYuwOenMdNH2UPiOWCbU47UF6
ZfB+++v/LOiBUmmG5qwxQvcCOqywkAyquseN2W/QUxfxFYTgrQzUuf2jYlbAirP9tXE7xCMQNWfS
I/VzW5IKNEOUCp2iOBWK7KD+PcKpgYay79/6L7ZDBV+fN3h6h+jseUAH2PHnOoEFwdbGtIOM6vAr
vdMVUdeASY6djgkLgJsY0gaBzXoxiX8H8MFxCmqAz9OB39wXzIvbVtB30JOYudR1IcLZ73GLEEU3
6nKC46D7omBGYKDk1+JGYwP6nnkLQbzyviqtum6T0be7USDu6atI+FfnDIqLEgwI8XZa5XqYMXMz
kQNCrJOiu63Fz+OdXZT0pjhwlztrH06vhMkx+tKSxe5RF1Zev+lpT1tkv6g3tkE+XNgROnEKXXoh
qYZCHnpsxQ7ZIBcnyny9zkk5mCF28LsTqdiaktoJoz5YMUEtCgRU5GPwks7S7KhbPGrxzHHL480A
NTcdRLEUfPhtJbqPeCCVOEMoHS54aagy1y8y3ldMhVf4i9WAdBJinSFchw9ZBRLtMwzLvili1/Sb
ac4oQ/pu4NPxZuaIE37hiEPZDL7j4CkcoYjKomlbfRQEXjGtYxmdUeD/V6//ZyOfqC4qy1NSEGgR
tScZ4A0HQbwm+X7uyv45Hh9NDVZ02pyjFK+i2jxsE8FO6U2Ukg00VYurW92gxRhiq3ezMXX81Wd1
w+SaqiwUWs1qckvPQW+P7NSfQAsQyA/swhrkxuhQMLNEbB8fl5BdD6DJEsZ3b4LTbR3kGWxK7ACf
T0oczbMHQwO4uC5tZ5rlY8iuWHSsK5OGfKjWXbLUhNnHjHyD4SjtT1ZTzKOkl0fMzZ9JVAifK4/7
Q/k2ZqGAYovYH614Yko7pm/+L4DW1XhreL2YaSaL5n2g0XtLi01kImQV32EMaCG/7xmdev8yroE6
eb9h1Y2X/d2Pwtfy2sJvaWEZW1aHil8Thf2HCc/mcfbTIeAGCLqQdFWTKS+lEtfSy68jwwQ3GiFi
DNhEMSljBuvMOCvdFfFQvPH+YF7f7EqOyCUrW5XfxHxyZYuI2/1ZZw0Jw0NStBD6yLHMrYp3Qx0W
dAY266lwmV6Sx1DR88InvMHl59JVxaCugrsgz9dVaQhYAW3yjREs6tnkYBwHe5bhMj5xF5RwUZUJ
nMORYn7t4FNypoyQStQVT3WLjigMdkzj1VrFxHcP2YSvVIUTOUSFLn9MEydJExaMAB/HJ0Uv1ez6
hXjAqyYyTuE8OGI9ed43YHhAcS18S3all6Bie2a4m5auioMylv/1tp2DxteCSCWMDREzqU5sy2jD
Ca+kuxofGkJ/fKMtx0tilWmrw/jPtOZbJy8ScBLs5icE3i+zcvJUFzlsEV5xdZZbs9jCtby1vPeC
/3pFADV/V63niiZUXUlGmgTh6qpZiOkVSR1qHEJ49+sOHP89IrYru5JjjUR33UbHVF9sSFo5011K
2MY2i+FkdPHakekU3f0U0bTJICsuE+lF+XEQdyjfx8ANZauBjIGdxr2fhg2bZ5zeBoA2UFqlQixP
FfpxeeSQaJJTBwc5nLA2gFvK8pnEmigwXvCJgcNZEtBS7wHWFQ6JGbAZ2I2bjg1jXUsEB/sw+83T
jN0LYi0rHPnGhBOwXIrmLZ6XQdtAipTe82NvvNOD0Iy459qm8PxPZOhJieveqSNfDp9rHNMS40P8
nLmGLTWmiqeihg13U7MRO1ZocPi31nRmXK85+HC3Kwz2bAlIbx/QSGTcLlJ3nyE5QRG6Jycx8FLk
0m/RQJRZAWs9SKx6GlpZh6DjntsRjoWXz4Y+Z0luEbg15lVQ/v0zqZD45IyAHqY2AItArnUgOEOZ
Fwcj0P5A823ovKbU564Lr69KpBx2ub/wirm7KQjaYp6b8eQm5Mx5DSEkEepiPONo6uslojwRx7aQ
bBGLNSVc2B8n9ziEpjMiOox1OoIWr5h5A0Nwf5Z98CtWYEf/1ag7W7ddCvPzZUxq2GQ7hTTED+Kh
jergDFsxkz+sUhUjQvEqe6RgdCbbxaz8JAscJtuO8G6sNo374yCUzKHS7R1h1EQ7lcmV7RW7iBxv
pJuQg+/rWcL9miBanjF5ZcU5F6e+qOiePaO3NV2b9CwXC+cWlciKjDF+hNu4Nt4yG/ZMilV9ERDw
RT1ecTNGDC220r8GQA15oRkKZ+NkClSBKd07fVBUejb4D5QnqJL0ep0ugsRoVDH+VY7gaWcP9IE+
WOzjNrEAhnSiYEZdwfktC2G6HuGtjbCgtyI8EDy2Pd5W8D1Rig7X80nvIR2TVezLHofYUrrfiTCZ
K0kZUq3/ZIUf+xYXe57oZHXyG1HIDX0f4tk1sqIeo8PvFeH1Z6E9mEXTFlbKzJ1sZMZJ4pE+bo8L
9CenTKvmbFTcHazuytz+6MAsirduGwdLYUseb18uuD7DjEtNSRNY1y8RmNBsbR/+wbkD6BLo6fTA
p26NS+PnMkm9+mkCI6uRf8wLM54ciiSvBxsbsZXRrKI/e0lGoBMW4zHXcfJapxTN5idZSC6PaLGE
dmb8kT06KbhrsEF6fJDbk34CXc1aypSFpzpThjwDRUWaub6kNbNcGyxSZUnZuUagl63oeTuVl3H6
VhhXL5uKBYRarqfZ7xeOV29+rWG82RMLiFI/vPh1ygxIF5Yg8v9iUhOT9bOECwB/okgdqNTCpZwz
R47luRtlbeCiUR5AUjsKp0+sidMc5aJzwUhBASFyws51qTMRVgqXAcd+jF28UsuRE8mzOq9jXvLp
TcKdOg2asBfQMlLCZRZv7+j8QSlAgaSFj+kzXLpZDek0SPxMePnezzRAY0fjWNMUX24ROB4IYjQs
iKmj9k8jG/j2zS3GP63fs7ufIaNopl16EpDK7J7cgKlJ8CRW9/hrrE5uwfVL6iqU+qoLdf+smCQL
K79QbGMU64pGFN8Q5drt18OCrtD4x96Xr4HFqVBVIWEloGIljTYmjNmoB/7cM0k5ZfL3tW2uxtAA
cIROo1GmuIQ9zNOQqGYjnforzAc3wJ9F3KZGh4dkFwYbMutjG9wltrETq8K29q2nE/FVAf4vjgXw
JDY8FIKfQ2lQOBeB8i/vAWVNlAqq+Qnb9jBduPp8gQi2OkX051P2FfpEsVRG0hNtJ5dznXoqVsLO
L+U7lgzkknV8B14ArzqpdXkO6jhn+lsba2yGVT4ZA5rNqSnqYIH34977pKYCH7XhBwrlnePv1CAq
HTBm9O2JahVBtWLTyjL2ABKvlOvSuY2rnG6cMuACh97nRPLKvZcRTk3kde9gGt7tR5Q4oWVetYS7
PBAINIZegojp0AnKMHPB0d0xpzO9vatU6LR91xZvrKEzDRPyyvZdVB/23eqEWpZjmXts8NU2Vza/
FbvHpAzNBZC5jnf89vVk0Vuo6lp+5L2f0w2VrzmtKUQg8S2SurJYWfoI7GyIIDZFG9ah0rVYNRKT
k7vjS84gNBj2C+V77fsloClwM2z1nuSJlBIfYEo2eWbeOLt/vTiul+/x4XP6yJ2jq3UAuPlgvHAR
gKcqqCg3hwL7Y04He71Zvn7AdcNpRUcPpB0d3gY9TdrRlTqSQdKXBPluAlUHMRaysHRE5F0tqiK4
PQZEnlIDZop00LL7nIs6VzwpRffBYGsVzB/liSKOiio2+7Ca25X0HwLldcIEDRziItg8UMmY7dVk
R48SXEz+khYqD0EuTNMADIa/FLiJVzoG+reKSOI5T1w73Ugg3ZEC6Y49V/kkHqDCbsT488TIi0eq
jg3P1bMWKox9pJSA03Jf1PeF16D2D5/MzhUYYqC7x0GVa1YKNj9E4+mWK4rBZ1ojB0kS6Y1du3Gb
O5Sp7pbw2F4Vp03H4GDelU02uccn1J4ctw5PCEWGrZYPyC/U7paC1/l7VM9OSV6l66GpNlaN3ZQd
vfK8Cy3Msm8EnVDDQEH9iPu6tJTZoe71tQtki0fpxc368I2dOmLU96+XygiE04b2FAkUVUMGOQfc
RGgzEPqP8TI2iyC02r670m6eKEvG4t+dX7oDBJ2Z8pVAAz3zN6wgWlgk93JO1nkUcJxkg2frtizy
/2OZyAe+pLYJtKazUHbY606PGoy5MlYiLr6uvXonYpsC4U71myAKYMwvbeHJfSodeoRaJbM35Ebf
+tv3iIeP7Z9F3l1WeonlyVibxbFZVDwctJfCT5gBxJMBKzxsSx0Iv9qxUH7GWlKgUBuFN3WpJgGD
+tv/BPyXpAcl8tjsZr7MDw59/6nttLIopnt+3pQF9UgR1ILVxoKxQS0tlw3H48JnrMRDzYJaMwqv
cZQHpWEVRq4LOYjbwN+HXSFXwqChrVZyv+4KgLZO82FOrcsdk6WhgFZ6PZREpmRlvEJLXnRP0rZy
lXyJ4jRPwlIVQE1waZIv7vlHrsUTpExamM+F9afXkSxezRjn/5LUgcdF0yDnaE4m/m1azPzx3UUJ
D2dhzvC8ve2xP8rKjj4VC1pSBQbGeqTQuRAh0gRhu/mDuHyY+anUadJywx7f7CxpuuyKb5MMq3JJ
iY3tg8NI7P8Bf7ZCHXpRAcGn/S5YYDa68gNuCDMUsBbbrw3Aknm568f0U0MF9qLJr1pmL2nPEZvr
k0cQyQkPIjUJD8uo49xTX12T8HyYwgYuDMcWVV0pGvC1A/IMz+3KDuJRq6cC0qhEOc67Jq3UAKYi
12UXnc3zt6C39rBgmHJs5Hprtsm/WyFg+IgIl12es5bzKdi3ysAHV22vQKXWRDJ47o9oiRvQ4va2
YAuIyb5zahiwP7jBmN1fFEI0E1G0HRoXp2x0R4Qpp8zGDKcrt0lZAqnSdj/XfCbNJJFYtGT68RYD
atvookkByvPk1YOvxLn7ra5VmxYRkYrYhoA9+7MR0OGgrKcQbHL3zAshUYVLZ8w4/Kk8PLj+JePW
jP8yu+EVJ0Z4Goa77l5o39jOjGsUCAfxu6X5nkoqOPYe3wfDdtEiyGqFa+ps7tv0u8FQ7jL0NcSS
zkD83YnsjGxIeTpQPIoPdMo/sp1bYUsqjwG31F4Yb9lBWPibIcUnsBj8m3C4RNsSxOCGkyVwdMoY
Nopj0Uuluxcwphh1agd4980WdNiFy5VkNgBwXm2DYNTDOzmT0IKl71GHFrgC3Bw+wlv9duUUxfA7
+9B4wcT70DsYbFE6FKMb/gsDjO1V+Nk1F+9me1wCCg+KL/OWJq5LvjUBHi6MYTYOziyEAmpe75ai
crVgRJsnq2ulk+a7TmjR4nw8U/nsNTz9O29DvVusMbb7+muBFXP9Ao+WdbTxfF1D+C6L61OzauX1
Y9WyQAvF/Cdc6yg28Y+VznuprbBY7S2/+fKNC3ghCmms/EHtmyskY50D5jHAJxqgMsTsybZAPOJd
jgNWWXascojRjMyjHzRE6k/MgsObKcx1cTKUvSZo7I2pTnLdu80bGoqNgbjuBhRZklb7T7NCNk16
SyQi6qUt3eiZYIZvcpQSl65F9qBuX65LtpvuZfmFnO19QdJtRNUat7JySOCP2CmlcW+Tt1BkvsTG
FPiNlYSORV7ixcg5N52WJvejTRo0vLXLrYo3Ly7Qw4ReFIo07TjVAEFJd8AOhkEpRyzDfCPjNQz4
vgDLm4f0frI45Dvk7RrWVfJJck2GyIoYN4ctVIhLVyyLvPCaWZK9J3JdxQVMSobojAi8qCwCyuQJ
MZkiyYtaanegqvKbHiD720+9fHitCSyJ8EQQiyzl4iZBKOxl/1INFH6wgL+/xnK7gL6+Rn8cF5lP
tB4grndE5KfS0PpoM+T+ViRAv0bwzJZMQGl5er8Puo905lw18yOZM4sh1tD/d4hdSxJcPyxfHeGx
hQGUhTM2HF2m3Rwdkb05guaxVSAWnwVGzQgQAhpGB2MrwoiYlh9iiZVkweSGEVaQTAwfMSta6yG5
QR+rC6OicD3XeStkX+OO0I7+oxb/RicqceuOW8oaduCl6cUZQi7uLqGI8ikVzsOjghxd2T2D5Zu/
Tidvf7dMtznbRddQF1zlZsME4hH/VNQ++XUWt10Rp35m3s46UoZ/cTv+GbL4uCI0Z2biuyp1VAgd
WzU/63ixoiM9cQ5hicV3pvaW4R6r985ELjBWC35OLcptFBFGjXHG4hgNWYzO6A7sN8IXQQKmaWV8
7MHiST7tNRVaJ72OVPbxusVbOS9GhtjskuCkbcXsM6yIYeofIz76TssUh3MYjAbxOpmPClVzpRKR
BTChinp1d5AXpc8O8QB7oc2MxC/w3IDcAumX2Y++6p5S3sf40uDei5VyRfKUpc/Ec1aExkenhw9z
a2dgn6wkLarkyXenkkc1MBgN7WHd8RBLTOCQgTBc8P4AiDhsmLP/wQoJa+xHci8nJ8Y8ZbfUPi/Z
XBRFrUz6cfSZDD2ZfNIOQydwr4RZTIdHqBFefPwuohQIsW3UvXn/Q0i8Rx94kwW+d5EP5YgcKyvs
kTH/dayXbEWHJYx1dLmLYzL/JOvF++/rzd8XHmsdJQBQOqnGnVMh0nZTJowuCj/W503g4eDuSAzc
RYRJe+qsBSjiuW0SEW6HuV8MgdWgmnC6eIdp90pe4quCdEM1ZDBFiA5l+2q4HO3hLrcaor/ruATT
IRQDeyzvZtLLgDCL6QVb3FD8AQZZXrlm2bX45uHVvSNNz+GPPPI7jARzT9enyorzWxwfwh/DHaTx
8RGO64/tML/O9MpVfOKLwwA8dvmVuRZuPQtWidPAy8ZCknMS1CrrcFQVk3Y5k8Q8PxraiOU3g9Ex
nNswpGPGv/wc7xAw08070tXUBLs94UWK1iEReY9sRyBA3hhbYzbQvXF/N3kwDHjVeQzdXVIhx1Og
BDif4X2iF6o/2Th+9M6lKs55Cb4AL4jkdNqgfBlh+n+3dizasL5XYyNf7t8d1HWX1zurd4Ra9l+P
CXcaJjy1TYSD/1vGoSdZvVnZYCVE4WOSXgUZYTyFVwkyGoY0BiW9Tvw+KmSvpyrfnEiYcg03iDrJ
xEhXuSX5rGvGXgXlpQ3lMHyGE0u/I5CPS2sSvGG1ihz8wHagiPV+Lq11fnT/bczAdLMDm7L2Uodv
DAG+RG9I0VLTPNCRREAn3OCFdW+LlRD2pHcKXFYFoMdFcTCkjSrIDDUkhwWnejGtiEKD+1Vg7FKW
Xnkns2j0O0/MGkL8NEjjny+m3Fi3HonAWcCaG7oicojx8EahstHCG0owzmGLWx/4gi3sTjLYD1ob
HPlNAolfzb+dkiIP3qj94iNYnlBwxURYsOMWrCRL+hX2rHBCDu8gJZX5hIp3knl3mgDp9uoKxDiA
I+ycw22N069HLfqC4mTvqMS952cyzefUHRjTJzeXNNlhgie8ENII9fZ/z3r4mjIn8TM5GwwhtwBO
YhTNPajJt4k5HTGx2/YbNEGKBpzGBhMp9ZXQdUY+oK48RJrVN/9Wj368U4PdnnVeHlaJquLK0EIo
VFBzBtyqwpBs603T42ehSC3c8q/kxYqj43GrZqLY5+mlMEusIfY+1ucrYZO2y6ssuJlzlMBPKsN5
3UkQ/uzA03/6OYJVvWhRnX5OAuOtZM4mGpmwSYQaUXzzHU63PH3OkDGBTPmJO7MNN9eVccFZh7HN
zgbvvIEp+rj1/ubAXOu1pRgv/iJh+OcBX7l/oPSElkVqcpw8a0b42JRsgBPdy/CQBUsizeyzveJU
+ioL/HgPKrTkAAY7RtM0nvURTP9N5hL6mlg9ptRvpM51MiSEl9TGyz6RWVBQ5D3wHBLUFifZZpnO
DTvrupHjiiki46Ek/Jmu3zXbbRq8qbzmWImlObGv2nu84n3GaA9BJj1bQGrOlZkGa4BS1Q6phIaJ
T3JvKn+IP3HheuHokHmamdyEExfGyk2TJlctigeUPyHCb2QAAh0cISm0/hg9T+LPUVxmjtlPNAMy
L2loeSPPm1mVppFRtebI0BbZXGoDUceBg6/saj0KQfpS+YDvVRY/e5L0C3LUcCK6AaRCRYAOfhoO
HOM+9/WBfWBa/wpOWyzS4zYCXY5FAhKjvnv5dbYBykNcKHebFqkT1+mmADEt//8Rw0jSvcXy/3Hj
qXnKjYCBo6FtP+UkF6FHXm++/SoMINQzp/v6E953c1dv6sdUlvkbzrpWBA/FY9kHDbJuo5CtxBDt
73B8ooWEnHiLLfr3iFcS+NV949J3ucgw1a2nJU+FQ99ruAstgZo3KERhqRkEwhAJO/x3lsAQUcAm
2pmcBT9Te1WAekWxAVhOQ6ROaVoNGln3L2hNcEQLPHbabaQqOaz38WE8HWomGcAKA58L9ZSzUNTI
Cs0lwnTvRXn4ZuOol5MeXVyXFcxbrcZUMLgmJ55DPHaOgwbxEAj3S9HPdFjJ2klPfuc0ykhYlK3F
0tS0YNE4iCwpUaqdVj0RVwhhCFnbvy/5dPkmj5QeHEs3etOqSyknIvJ2iDoI8JOrOXPPhVZq8wWS
F6r/qyCvL2hMN4KhkEoeCSQrO/mCV41LCS/PqLTi+QM7nJAyOZqp/fAYa6xXzTwEwGg8v2zTsx0w
5fPB2btYCaAL4FwVepUrujnbcM3V05cA5cIXuL92+QvOVpU1BlUaWPCR9NjRuz6KMirpRGcTv371
hO7wGTpqiKhKPLjOfpjiCIWI0XyajZ09lF1Q0XRaFzdCs8ZH0/7kmzc9FIzHu1C2GX8ZIdm5urZr
4ED0vhiLGOWQRxYFEDOjQEni/p6uY94R0ceXb1pOzzB8Yp/CBkymXzeqnb+mlrC0EX06I9aUKjhp
PJEk8Cds9/JiO1CPnA1i1bT0jcS+pvI+qYurwUU+X4Dc81Tv1RNlYAdUkA+Mu9vSTg64357gyVZP
UkPyexeYggvh5upv6GA9vzb6oaaKWw1f8RWNlzM7hFBv7Rbrvql76Dy/X0kAvT4o11BKiRjr6FMj
6o05iM8Fg1IkPGHp/oYylnfZDK6uF+jV254uPOABA61R8CgAvl5VXLpoyKd+zQkotav6vQe8Xs/N
9m6to5MDuASUB4oZgtAAysFMrHKWABTV8fmnp0WWgysQDH07nPV5OuWuRRsRmIE0ZuKCj9FMzlqU
g9/iH16MiqN3kBxRDzL98/5dmDk096KE6eGX5QJsr2ZbhPtos8fotQm9DoKLQ24Jjb+vFUW0RHmK
uSFfk61bbGqkcygkivSNozmNRbhvcNkZeVWk00otc4mnbKOHeihJOspoXxm2nmEqOi8vmvyxKqLi
QIxArwd5m+GSxxBlbP970nVYaDCZP6OA1F/U1XQ4xDpSqJRGre18jdMPhgLLHBptHv9PjiJhOgoV
dv99FAg1EMFlOllPxzd/yFtIlGbQAdKqCkUlSG2yN8wRKKiSPL6KXSLV7/9tskFsT2asjYj788bU
6K3v2vgljmyGtRPmqomv3W1kNs5EQXIhmQDfUebzoXXvUZ+nw7FiYvwC//Em5C/ec/Oj+AQq9XoB
x5jz0faybBatsvbJxetQe4lyWuSiQbIKO2Fp/qP3L+sSEEW7V6jTW+h38M9qpVRgPACxfjWmUXPg
Q8dS1yZCm2FiVlK8TV1xN36gL3rEHevT1/0JWnMuaVbD6UfCYotjcNFrADFnrFCUoZBEeve7wiDK
RMXACdKPcf6vCFRqCJMqwyacthpjEmoaWVs7w2sutqeQJMmb8cxciJ2vfylwAGsQxZm5Q8cpd0yO
LjCTt3kuyKFngNJC7gxA506qo+wFo+aRXJQ2b8l3PXoauDBVpAHxDqCh7fvxHAQhe8vpKo+t2b4b
fBKp1xJpus8Y1eoc27Z29l6vyTrvAbMA2eSaFNVZGOtpQEC6vqWZkC62DtI2b6tYmZJXMfVRcnW3
wCWqMBJJLqRqtXg8s+g+9gSw9DpLxbOLHmkvWqqlONt/EMCI2Vs2NCS7YRB0BWI75gXx3pQ8BPXq
0iImL6stA4RzHfkGM/HUQypH5kxdKWSXGTCsyUUTRXoJREQ4MQ5hStovhi2bUsWVHj98l+4HqJp4
WRnXRA1ZKdTolWGQNKsyzXx9e5Qb1O+hh0Is6UKdtJXbCVTuuC1H5cMwTt9rawQ2abOXs8kluGTE
CDeFVo1nX/5bB26X0uQBK38rJjFza7HVQHTOrTBJLXN8j5L86tsMMv1Px9p/1LLpXEuqxHDQJzAK
zmwjryitex3zRBEvDYf7r8VLxPOhSGkk07o/eG0NjqM33Q6q2o94HvS5BxNVrkJ3bOPxKeE5QelT
TBIvXaRzBPbC6NE/twfYSCTCGamXkpSESREHl6VyPjc5lfr5CejeZ6pSgZS0NDtQkC0uRXNjDTQH
mOwR9HzDKXgILFxyx0MK6fNj983E80vHgD/kUT0Cw0hIThm4p4VndifYevuDzi5YZPDRH/vaYuSo
7W74KboBlE5ecwmS9BtNk/IVpAh356nnjr0xupCV5Nw1wi7bP7KhOgENPyXNCCz2SOvxP3ThyiOj
l644PbYwEzsm0fJaIBFChbRy3IDlpwi7uLzoyXw7W70AMzMTLf4UGNCW69Mw/93Ng5+YIxGaBEd7
ZWiXBFaRpc9k+Ah4ISY+ig+6ohclR5+UdT486gdJAvfLo8T7LUMJRUjxpHSIOXVp06UKQyVbd2GX
BROI2jD5n+wfwPhRVh8FvyYnwAqp20b0PnK6WlyQqHSzsOXUilvLpeRqutPxGJRmwBew18voS3Lg
f9X6IdCsEN/0VmwRdxcx1nfETkUYEfYp770WJIInwU25SClGnKilMFqlRFX/N8gVBk811mWiv9Ii
qj8hRK1QtanmGZ1Zj56Vlkm6rkpPlSX8+83k5tU+Pv7zzTbP9dt3pOig6Wmqd/A9/dczL+Ji/5Vr
B3UALLp2TvSZpma83qaJG/4HLlgyb38OpDrKsIRDvcwAdAg2pMR5KgBsdTgDpJBhLVIudJ+TKfH2
E1RETmXHeZmcJBFZlGD1hLA6UE2g748xSHkKiXKR4Qoda8X4qFaiirvJXUNkJqXM3RBk24U/4UZt
wfLvYO+/DCXN8cA9a4UqCzyN0iej/Pwp8wPLt+UAwkAXCNLepBNyKSNKzbep5CbWQvGoX69GuRPH
QYQtTgFXKS31GFhAlehSsJPnLUi1a2o4+WpGT4OG+INGw4x2D7Gwf8UQAwZMvFjZXcQftvH5/8DJ
hVwT0m9fuCpD+YBIguXab8meNDlf0Y7Gj6sU8rtnVlMivyq8oKdxzEIz9DNjPa6RnYKmKzKJiG2j
o7MbjB9Fb2YVuuiLY/p1onIwzKAHilbPNAWbcc6rvjJwJwa2Z+IGC0AoeSDlLl45HDRLbfDW1413
ekWjr47RZuAppwyNFLhSL/+mDk2wcz3fOV4oZpEFZifnhdZqkQHwoN0gIYuJXfQQzjFkE5+zTlEU
QG0ZUKWXdrHf1T7C74SSTrpHV6ilgkWt/pjpXrr9YEpegn8Tvlvirn+cqxarJUwqe/WJ0fuOx8yT
X9LYIWaJzCvsfjQejLjehcfetwq+DR3hUb5+XDqi+qDHZtCWPUHPUnSaapWUD4bcIhSMal4ifOdc
/i6omo9q3lKT9Kq/E6stQkvLJCCx3KjntOPcfC2FfOfZo39sBnjnXIOxIvO0my1Gta3cK0N7FtIW
MfciV7tItN2Hdj7OCLDPWDQHe3QgE+mmeVmXFCewOhuQSBXXK/LEJcS3AHpPldard/YUQA2ZSR+5
XNkF+LH4yiyRR5L749MzhL0yKB6phacVFaTP5ZDcAUNg5OBBJYbmVXEl0ux9/V+irCwPHbNt4nTg
IBO1Aud3DxX1rbDYczZrPUj0UZg9hHJnKHV8Gs8pv/7dK/6GZEjikvpX9074bN1t53c06fJL4CTY
5ZhyJhK5DTI4vGoPiZdKWeRe+RJEL75hG+52tg6M1vdP0znLn7LfLOjNIops0mYZnun9DHNz/rUn
fSE/39aWrKuBxBA01A3c3WQnRAek0G/VRQO3lydwbVz+h68C06pQAj5UoM0PVpHbjF7AuA4EIl5X
3rPqDHgQoluxgmpl5CnMz8qRxJzJRQF/o59x8ujIPzGrYn+4LrnlYzVVvILF4/j4a6IuOlOYW0UV
1Oo0uzM9vTD55OVfsdLBDTAnnYEscVqMOtIsQYCwou7Rjfdstq5meL61tw5Kwiih7qbmox7uJwgk
so1IVJqGSiUiXfZKl4f9PbncOj7dcwzX4I+k+tc8pYz95cPNzM/TryljRfbmqkL2Fc/bupB8cScx
Nj2ONi7WO4STXJWrYswxMk+3c6k2/yNFM9S7zfYxpQ8lwcE6wxMMSuq8ByO2sQng5fIvBLLPzDa0
hmX+kRkO9/J4XELAzfbBRh2Pjp94nMKMBVSBphKZKc0XZo6Jy0ZpDYNNd9PX6GhBARqMcK6hiCnV
d4atQO7wV5rY4NWcPSuuJrSwQ/QlVrqLtYk5tjQYRWArnLFlqZeRL/u4Pp9Rnv0Qzd4dk9/tNwXb
rlrHGe53M6nOKjct3Q+p6pbxJDLvZehyd2/u+bzOAx0+k0n7PYCgAfFRCRQjax5VxW5BIwFNg3ln
alBtfDTVWWhNq+EneTAqUkv036dHqnV0+apgXfMwQCnRE757bktNLTXKn9Hw0R7jUzfHkGWfCUG8
Z0El3ul9pP5581ODGaXyY+ioJD1f6li1gg/ro61oKj3HFbYzA3mYO7FgUxJbLuaH0h9V7BbJXMQN
FerjeXl/WorOHrSqbI5wZcR17J08kbwQfJQ1oWv9AUqEWlpqwUVjweWydqcSMYQG+K1G8NbMM0X5
f5yzX3Szteba/l58RdGe7sEa3zjhSbxfZAW16j03sLwm+vfo4eNDtMjqrPlxlVxUSxpLs12fqP3Z
0caMDq9a35ullHt+Yi2lprDirJpkvv8zDNm7pdQqcHNaijTsDX04/xEIvq4fSwWk85JxOkxyfZ2w
47Dzmij6WNWxfcxXT2YYUIGPgxXwqV0QvPrbIpSvZInZnZdNKFv5R9iGFOV1r8CsFCw09EIEeAhi
C0ChraOCaBEqc1sdL8C3/scGck43avxboA4O7Hf7tPmkiha3Pi+pGPdDmpgIOPrYZi7epJWN3eDj
DYQuYwCpoCOYJP7DdT+HIbiqDJJtUWKJAbbdj1wrE6Y54unwoP3SqZ220k4FDXbEWgBNAdL4t84p
w3O2+kVHIHs+zXLTL1OUlF7mfF/nxlC4rz3ZEQ6TNHTC1C1i4sUoGDCJQQyN2Hyeu1COKl6wXbY3
qj/1KZ3+fgUP32nf+A/rwoZVBGARnc3pzZGdmXGZtza67zmjwq4m5/guijlVHiTLYWS8pRTkUNcN
s79P3AQmMF4mhUPY5EbL/drVvCsw+dbIMGM4Ajg90z1TKLrFR+JnYrNMBEWuZ8U8Lky81+LKCOWm
QciucqnBlpDPF5UbsMCHBth6inbRXavbClQthVXSIjmliqhUcBAZBnTbx1tlc4gpJUWXPrwvbmOz
jziAZTu9xcxbE8BKAc6SoEJi/9h0MeYgyxzeLL6R6GJtIwOXNAfIsW/7phs6GtPqZ5hyMUOnf7pp
vQw7IZ/uXzZ4Nd7wDcaim2JQ9upwOkt3WEchHpWcOpulFxvXq7ZkwBawJ2wf9TU2vxkCZv2O+bDk
I8lE4v1G474gd5tuSIH4D9XZQoj+Nrww+SGK/FAU2q/U6RrBHhR38UdEibbXMFwjQBmnz+RM7J9/
AIokHlClfG0BMiGmHtjwKaIHy+mjAz5zpeaF0AZ6YORp7fj0yuzCyrD8TjMntyw/4iXyf8d/q8N3
XHbNn1NtnjJB2Bh3hZFJkPcbg97iIWAaO5P8ck3csG9l431PSz5P2UMlT0J5z8anCsncHwQTQshi
yQyrPobJMpXmehgcAYkeeT/5JdXWO0SBa+02fpr+055V6mijrMWKp6hBr8Lm1Es9vgWkWbx1Oj5C
n3nL/+dXfNTEsAoWXWstNmuEGzjfU5V7K5O+3RISRTGNIcq2As9WttaDmJvGSKj8p4siS3JXFxiM
RuFcIUwkRumEfiNaI8In75dFOpqg2a1zUBbJkGV94vwcE8eckTiVzM8bhoUekvpV6iEe/M1Y0k3n
JjAQC8wha8rDtFp2YzqyHl3JeaOLuTYHywiucJpmoBYo/T4dYs2iQR1AywCEDcakSbWSLsIQm+2m
Oir+FyMW4TK+idPCWNtmMNtHTDHGhv0BhJvhEZApcsyTs/SednjEhCWB3+lTVMNDYxM9A24W1mJy
HMjglTbSyw1akZ0iE2InXxd7bMfhcsFc+d8IC+zy9maP7Gm+Z/c26q//IROYyZp7bVJNG355YLFZ
YvlVqu8bkaFVPwkdAW3oCrte7A/1RLfXk4Lp1cr9z7IHkbFgqHYyO/jNznGZN2v+t/Q5U/FQKzIi
LfltHEtZ4Bjhc2DZ9gLui1Kev32mheVwDk82o0/UOXYjhnGTTf46cO/BIjjYa/q9Mrhp/0vvTnFk
A8RaFIMwjdV/Jeu+jMFe9SCRVyw4UbjDqurDnZJEC4s0R80NvAWBveKHYM5fpk1Za/KI0ocJgZ7j
ae3TJqmu2y8BV2Gn8h47OSNiOxtSORbfEDln5pHYTUlsF3Pz9/roaPONankmcQiATRHk0g8e7QKf
g/EHS4O8qda+MY58TLWwrHGYUg5VVwKf1zqmsFWDFO2DkZ/08hxFl6l+EbomlRcnq8msXbBdwIU7
mXjTZZQzyC9RLLwzp9zJtZiOeO1R1A/HiWmCHhWjujnnGtuj71k8PwRedes3gTOh5Dsl2jwt56DE
qLXFHwYDcm+EN6m4yuehhFZam4dJZeA+8xb3PZPukWWQoyah7EuE6JhOz4lAED1D5QNrbeLbb2Uh
e2Vbjrge/RJIgpq9csM8iXLzTGbLaauURthLlQCDCVv3iVmyCTQAESmi/RWsKB/w/8QFHtTb4YLm
qKa9FA9tFyVP/Nl6Rp5mTrAuaJjA+DnERN9h/6801ZeO1pxzU3Tpul8PT5/z2Zzk92MoUOYvMy9E
EumHElG/hAvkdbiTi8tXdmTXkS91qrQd8CDp8JCD0yy5v1DqwOazKE/Jf+ddNa+BpKq0Bv7kVRZR
i+sEoAwMnEV6/IEh70cI4XgBi/EcTETKGEjKC32ikSulcI/2iHZQ4yiUwZurCMxYAPfjX4B5G2pI
HTkPySoUHnixS45vsrKaSUhd6K/kYpHuMKLYwsIyyYu/lXlUcrlQzv4cd5gB1yJ9pDiwtXBluydx
LVvisdNjNEETWLPDzmBbWM2ESD4m0AmBgYgrcqCpWjZagMf5qaItjVejxvNmYzIosZfvYNWR7G45
cQ+lWFOMSDogzZBBN828roIg+IuSIiFQQQs3q1cZjDA6qHWYvQiEA5WfR+EU9FlS8m9g1/WSHIPe
PXZLkyeGTgF7jabTPv0YFneFGfj/UoNGy71K83QBkUTZtdondV9mR0UrrLheBAEYIh9Hx84Qv9ER
9NnLip5uVsEOTCcLzrHymZLqiVQNbo6dPIL6KA1C0sr1tERDQclIovBAQ6UzSkhGr3BQEbr3W7sN
PBEWgnERSLYaI9Gb6VM52Naa9HIwtBV1LtyeGcfGwMWJG35JHc5vYY5Od8xHDRxtEusHmcUd2y6Q
I1tiGWrlpxbXiGD3FEYzwQteqASYceHroQC72dzrFQmniu8KvWW7XKdAqtQea5QPHe7k0fP9TWEt
FJNZ/oyoxP/fENglL9EQxSDDNQVVG5uFxgzoj0gHpPpGFROrGOv3FhXO/5Gg6/eIIrQZLAVWgDyN
cKy0L06ukTCRV6XxzOoDlcj/uRDUfX1OIG7dlyc4IC5QvS2ZULcwqIYabxX3NIsPrmd/CIhZXvFo
2sS3BuJwsk1jomupJbcbiVtfJqYkHzWBjp/nx5Dxu5NDLL/o/ODP0lxZ6Cbz5HkUYOK+mfo7Hk0j
WWIDpEHYap02uu0oXkJKgHByqkuP/1Z98Vw77fsAY0XRNhQtUKyWoAf8h5in7RC/jlSUQJQZhjeg
UaXa5rKB1dZhRbHybGImSXPlUzbrzNbe+ilCXQ/VaMoixw3JL/xiF9XK7I+eek6blj/g2v+EacQc
bEAKsaMbFCu9iEIUpeoqKudt/IaJ8yLq7qCgcKwizSmm+jiNS+LkY7b0+Q9Hib6h+7rQGsTvOsQX
hZPgWGHTAJ3Af3rsv2NfnJpwL3Ul1iV0QpAvzcpRAI+BIS6varR7XkPakD0hZPoom7uGSS9XL++L
xjevFjnn9z+7MROFruVyI7zXX5qDzzQp+Si/wfxa0tLhntAfhj9yhhpelB0viPKMnNQp0p4errFD
Xbll0PO3k5xstCmohbpvVxYdMkMjzahKHWVIVBNV97cMaLjpzrw4ZUPh5Bpna3MvkKGEsEo58U1m
ohS+dbL3lmMeHYGeaj3vanLa8il6NaU0sML2JRDTU9rCletJtiEOafGn6x4t1pNh259LhG4Wyo46
19jJjy+MnUFxUjrgfCpp92an3L6iUBTLJI5EUN+9dyjfO6TCwgYJCCz/pJFWdV52EIazvwT3kKgo
WbV9LN81sci4jcfXEp1fj7PmQ8zroPy7UlQm306CnDNqrtFdP5OKDEmgUvW6hRYXjOd6meAJYZ9J
8IDC1QxLuPHOwXibyofSnuHkAiDiyp6wGiRfKhE61odHDTvfrBTICY9lzYWynsLwwM71Wk9kzOtI
bupQ4VN9v4f1lVRVxH9rj3QexyvafUuqvV5cQqG1DEDlh/Gld2N3Fz5QX56oUr5D/oSrV/EbRknr
q/8DFWQY4uMH+2brKh5aY3hkaB1TCBBChnvQXGtDrcKKnNlTElSAeaR8WKKRGx4iPpC+W61wL1ZN
DvJkNmgw3ZGwOawsDG16VMCWQ48ZkS2opUR91jO8dED1oHXbcrt86t5t0ISEHo2jUB93rTDKbvuN
u4GIcAtFJ+BMranQirU2eRnnTu321epuTZO1oIqQdHAHix4+0Rs4lM6ao2oKyswLQSqD1bUh6aj/
hLkKk0Jxhoe18ZQK+Qw/eEI6M2NOFLW6qxAzXqqnl5ToNaWug9YxX0FCN/JSvnhnPOvJ3b2uTps3
V3ae/6s+RvXFUrH9LSG8ZbOPTynAEfMYnBsW+SukgNqrmuxBjlua8xXpWla0cpV5vQRU4NclKNF6
U6T3rwD4y7ZH4/xuJf/iTnR3DF5T4QrSaKGubA/nHjewC6t9/6gQU2M3Hn8ppTbS7br1oobRfVA+
wkc62srNKppk2cxODlXUF1M1YxO1UJ3Zc/6NIcPdc0R+bVbck69TZRUf6pVXX+xpdc1D4RR3GuOf
pslVWBUA/d2JRkavH3JfTr90O76rvN5USe2TIha5J4ivEZzTBiafsyHSTKrur92gjqIIzQQGKp9A
FPcALssP4vUZaqC4lHRDpRn+56cwzJOvFVTNplVh8cJ6cMQcNogI/0R4Xhv0CWcdRTFYnls+TG2M
vM8IdfSd0xKsG6hW+xtJXuEQ472Bo9ySfDGTrDWcbD1kqtNMfgvcrtnFnU/40pRa6iHeh1gt3KW8
8CmNCqyuJN6OasBsheT3eMwGHDCuZ5mL21nyO5pGQI0hZABXXwq0hNWPQbAjf5GTOxzvoNb5Ki1k
wNMORdzeK42TmIQupGxB27ZyzQz85a1vrTZvwNJGcfx9cU/9FlSIdDdCQBtVZz461/i0T1Wt6smh
6Bt5XbZEAcxEIY475WK5LvRs9i0axlOklGs5T5N1S/qaIdwxt7XOPVJaljLQ97z7MsWo8ZUaAHo+
R/ZZM9TZzyEhJiXWjZzGEbNyvFYkUAuJuL1zpLgEkvXA3JBlEvnrqKMN2/Bbn0ifurbwVJq7+t/t
dgrgQp5oLbuujhePjCGnNUe0hIFZMqMxy6NsbcV3GpXqfDR4zZa/sNTMp5FBYR6WPbpBqBA61B6b
H41+us5+can9qfv5LKJxDRHBFksRtGhP2UCi8UkPkfE9HZTsgi+DPaNsN9dvIJXYAnwgSQ0uKMG2
mcmGfdAld39hxyq4+K0fyKFU5wt8swlrA2qMDYPEtlDAIH6ZTwZ6Mq4sfN1WXyv04NSgL/KZfoeu
7XIDTc7v7MK0CQeBRxmws6CSbtM7ZrG8Ejz4N1IHdpep3xtM66RpmT45ANZMzF5gfJl5/cepnyI4
yyTLO2qeIaTzJkd0QCnoG3ggQPGKaGf41w0kaOMZfdejcavLWoduAFm9qMIhRIWvNAlul1FH1c9w
s1GSY/Op/a6ywGvJLIkrjf+Ty9a+SFqUWe63WIpxRARGEVHE8lTbYsWopA4vEKR+KWwtzFAulJUi
P7cpb65SSBAFbzGUzFAnIeiNxxuC7hiNPCRnKl8F3hkhgEMgd0SvQcZZ2z7SfKld90yPxFJbh8f6
g6ub7b2bs7s04QWf7O3nL6jeug5QvZtiL0go+O9OWxl/IC9oB8forjYvPt/0VxqnPAn0q7GvYmdY
/VSD8aA/qsdcl6y+uIA18SDp8/EGx+a/f8vxmFa7A4wFagVrLovQBGIQnhzUdSbK1mcI3txby6ko
d8DiO0+WnLYlEMWyszZ309m2nEAzi9whvBuRMpUUr3/z5ntGCxr0X7lZVdT9VhCD90iS82P1qHpQ
GsZqQbKKNU9A0x4FWIoHflCat1aMkP3K/rVXLiGLP1eZz80UzaGcw3io11EexWS914i8da3hTMT2
Pcu56F1CsT778XCHWPfTO5N4el2LUg/VjSqD6m6YjW/nXX7hAGJfkRn0jWQEWUXoOL9wCWaxw+8Q
yDxVE9tSGl+zT5mmzOZ6w8IHsdaLlDUlecaSkYsxbIwOVdY1Mn4OiBCBAr83f7en3kYPmziuj9Ak
dV2MuhPsKeryYvVdUrzD8xNth9xJOv28y4Xw4jPPEj+uP7wB1wGTuz1mxmYxVbXdcYCgcpnet6G2
+AVCRW20ifPyY5U4hYK0CIie4kGBliZmhnKsiwFxB+1arXkUg3FPypnWMofq4OpCrcCxgqdlyQ0r
j0sYSYA91eSJIeEYQgSY3r9g2ccUZOLtL1HWdTXFzgd8b2yIdRjhZ5Hja+7OqFEe8SYOKssKXuPK
i2WGjPGXs36kmhevtiumN7mjrc2ZtKGenildNNRDQfH9nycmrUsJqjSiYokxfXEedrrpU0jEnp63
pI5iLBjMYBELWuHvXHBReQgcSVKiMipmexqIenDrpd0ndjzYgauOI2HanbBROsPwhPkFcu1MWCcq
GS/1WqrfwPQ2Mt2L+60nMIqQFZQUuzPksbxedAeEHMPrA1WGtDYULsShGRxqTQeg0nWkUWCRTW0h
Bbg0seztPHO5FljqTweEzC5BPcnSV7msnUJos9OOe32SDRcMtmvOOzqqp0PIGvQk/OxugtwTEunR
uZC2EH0PvkXGqaO5eu6HI8Uw+1qickcVX0mn1MdUHJEYr/DjZhjRFWhYEKLgAOJWyhkpubucIFua
/YaaiXAyygMYv9mf3Y8rifaDYyBpIQoTBaEwYNhbdfYPZo431FgPQqh5q9YXxWSRAK1WJSULT/z/
kci6WlMHPkaVfcvfLOxa5f5aTphMo2c31MbuWoS6bOJQbGLGTv/VCmI1cNRBsTWIDgnZKlcBQK5Y
8QcVim3xLpb+ky6zDViWKdtTyJeTG3IUFUxwECLX3vlS6dSq28BnbuPN5/+YjLSFoFWriP4wsw3b
U1FYflOpYgOzp3xOtSjptdnszE6m+WVVu82v9EJa9JRnPYDqGMaLwLxZuY7o2M9o5KxLMQxHFQQK
vWEGUE1nVZRpFC5QAwYczBxXXoljq7LeF3PwoeFKH8r6Esgxq3vXnphbEgoVkKMb8Y3HSdUPTd2L
rAFxSDYv+aoyXUxBBfyQuyRekpH1XfbkdnLcmP/tRhx5aIgeFmB+UVVwqb/oAQSWqzubc/++Ei0T
xg6ESQd75L2jlKkZxPQGE2kZKGPnZG3ourxk2oFkWUnaXGkew21tsw4VDfWswIfy3nnb1pd/Okdi
pNsl/1EwlEbHh+eLVBtI+Yv4RrkbwSh10UKM5AXe5nGkjRFImLsWtbGtWAjipOwJgdivoDFIUuK9
NuWr403OuZHj/X/ymgTXfVwpv3/OeABO6DGwInTDNi79KiuLlOGO80+ZbJZ9czpTFWGZAFqqPjcB
rj4vMjlXE08p4djl8CQeGUC1XzEpDSelb7EFiAma2GU+LKvI6Zd+IsEieiP1uY3eftNFwzvQ9rsH
cPkAbn41Wxx0p4/y+RRnR61yW9mflDiyhRiSnjX24IMZaiKghV7dGLd0hCdBHd9EXiIb66tErGNY
jciUnb1jaAzgdv9FD0hPE6xUS03CXXqto4B7Zizf6p8TEMNLpA62h4mwODYi28L8fGzZHN4s09N4
eF6SffMXVWFzZSLpIspopY+tFaQcZlfNjN+BUWoPcJjOpdEEy6HlXO/LtUDdsfAfItXhJzeUWuIO
vbNTY+SBnHNCG9TPoTD853RCma9/BJ5CDJ1xYdd1zya6f5h+b8b6gnNX5E30xCBRg7hicNRu3jrQ
W8w1cK89YQf3yldGnllvHDiK7F9AnIKKRspjsVJCu6zasX9No1I4glW1+9kUVYRnA684hQ1El8p0
f3Ge1eixY/PCzOSuvIYZg9lUM3nMxTTofAMu4dGYprV4IZotpUZ8ut+4UNwWStZNWERwBEM9RVFl
79BpGsdQZGIwMCPVVLi042JKdFySTwYysTlmMmyyJ7TojwysijoSG1OcFZhGKdWaBpPxEjFGvzAh
YgACqFFlO2fqU/TUwhNsoSPCFAcIhaXaS77LACIRzcNgFfoI6JKxlyTx10WWqEpDBQyJgJ1i9tY6
HmZ6Mjr9Pi7heuorgNov5Igtma9kh/BvE8S9bPH4vGDu8/oAcrG+6jDdvG6YosPAYB4Exb3/VnrI
RmtTaE3QM8A9ho+1prffQGGX//p+gYM7ESqUpGnQ3FGyg+CZPxYRgRvXTQq5HfE5JVVVtmCusTh4
2INGK8ePNXcxmCN/0pWg4WFwleSTihL1miJXQqsaBNvRekkodbISAXsLSjIHJGiAf433Pmhokeet
ru+XXoD+R7pNqzrOvVwM0PSxx82Hj2SAys5hEThi9rBdck8Gc7ne7vem1erZtd/BGPE8XGAXb70P
CO3e6RmYvLmOOCxNzgw9cGKEFfddW/RzkrXdt+U4FMDAl03ST3TMl2m48pnnhCobHfS3zibCIb4k
wBi9IXQIMHDb4Z3MOeHm0aFzLni69ku8mVsgy7EVYV01YOgpmP7h0eQR9F4VIRtR5xxOZS8Wh3LS
R3JbvByUz2Wq1INhTsxed6qrzk6hEtj/KYGKcqACGkeOKKIrqH47CswZgbHqI2P/8GYRF6T73bnV
BSMch234q9ZGufc6pwVVuOEPOB7WJZgBf9FZumNEeagNFds5x47DmTQA0t1h1bZMYcPa0t2xm9gD
dFipvUUqEKRTYWlJdNSR8Lj+kF1ASo1CH9N5mxmOhWLIeepo8uk/H5nWwYKtunLkOC84g2BNxfjM
TSGOkTLTNL3ljhkGSDlAkgarmHcH9PHCSbcRvC0HGJXGD8yd7Z/ARWAA443wCVpUlq9Hk/z9BeWO
lnRJOEBDHumkI9HNmASxZjoeMY790jNTaP5agt1H9ViAmFWaX9LbhI7Tp1iYy4HtUFtL4NzJI9Tn
R0cFmWAbT8yNGVy2pWrniD8g2nqcpK901qIfpItQ/4RFEhYMXcAynNKtvtUwFYbDDYgzGUXafKt6
qsmtWoKpplUETZD7Fjs2K9lNQK7lKh68GmeW/V/f3BW0oUqKYGruh0heXBWh35Aifka8y+2BSafy
MHcfUsXgnxf28+SyjKDtOyf7qyppf/yua5wkfJeVb4zAKejsqe61xrCEErXTl13EAs0oAGt8F5LZ
6daEYZPwOlzwPREM3Apb4GQ+fwcZ+rvULj/oPFrnwXuV6vDwP+XNTlFQaOLjstJ6HXIxb4Wh9Auh
DUhEBp1l+gSwJ8+lUnUH7sHOgA4E/6811fhv/xDPkgMrSRK1VJNZcDHaHdK3EzYhL3QnDVD6fuOO
C4rJqkfV2pvlbJ+9uLTG11O7vLYC9FcQVYrdkBdtRtHEt+RHmjFM6hvF7WQxQeI/qNgI7lNlacSd
2YsD1DcaIngf5zEkEvJ3M6Sm/xDpWdCLP8S+l2mTq5Df3aWo7R4kRUNcbMy0jipAeT93jnhYmEL9
ujwJxmpX4acgdY0/5btnPcYD5z5nI1ih3ijQsmW4/HaXxjb9jLG6py1bzX8UtrgxaMB/9Bho0tHy
/VB1wmmhKlBmTmtsTQ2YXAb4v3zo6YmorrrN+F2IQY1NYwhGhnhf8ij4E06xpMdCxh5ChIy8xchu
RdJJhN0IO7UoggTUBw1P5TGZSyHh9ZSJRFUsG4o5KZSzefs/JBgXHs3EWP1kGWV5Oku2L6QII+sA
Q5WhBfTh/AnZ5n5QR3OQJqgu+PWLYNoE3WAhHW+3EfdHVvl8HZf8WOAL/+giQO699Z5UWJFYJ9U9
MsP8WHkISXlnFxGHH/hejbLAN7rmtoLUmOS1pPOJtSnRLNdGkwDzlazAPANwEPWPekShl43KCu+/
Fb5Rg2BoRhoAHJAjD8ZmLxbPvXhLEkO0sNmn36jRqzNq9dneuDuuHfM3446Fw/p96MEksG997nwp
CusTcT6KkFSz7/WBRbxzb4atiH1vi4CgimMjjyERyFn3PShe/NnaqrvNADirMVvEr/CLZ97KFOxf
6WC1hu4P30OBQAusFZSa4QzvrNjzXTnNAAb5O0RzBWiggnO3ijEq8hq5fsohxyyOle+YZx8vsoyU
kaCm7z+CQw9+jTSz14mmLAqP3V47Fydpwnau9upv0Du4yc+rbk+AkadGDiekAa9c7JQlLNkyUztv
bo6rUqYYlb3PAruGRaqX6KPo+tpds41SopB2+WoOM3QtXMtK2x+M7eWU0+AFi8kLFcRiWSbe9exm
fTNn+nz/wUu9/Q4SZpFTEhXxtHRo19FBECRUSjlHM2RNjBL0qV2NcLRmPhOQYQwPInbnK8deHCug
uVicRc0ulk7veG0FSx3e5nGuYj3ga7JoEh00EM0OKFoJBoGzXtPWbKhtYu82zqRA0LYUgS4xf4l1
K4idupwcgoE9+rinoc7mB2jBSp5qy39iNn5wML04hFKEFSz3e5lHI3NEpXixetZbCC+8grcVY1M5
RttReuCOtjzVR8VnYXLYDHcSOHbjR1KwJkZqQJtUebeGzly69wAAT+WRO0p+6u3v5oM+izq7drKA
f2LRuMT6Vk86ZzVYK05tiVsQnB6tarTI5DCBhAruTnxyXrDhOwKjeRkwphhZIRhm25GilqUMSQWj
hp/nBiY6PEvXUHH7H5nHUhvUjjCRU1GIACS/ki56ahPtC0msjKsQZ5JB19f0y4XnFDRzVHdQM8Gc
8tsOMyXrlf2TEqEnKGWKiYbeEiwbbPpg+ssKmqsmP6Z4t55o+1uZwNGkw6pfV0XkvE1IVIkFm+Ih
pwJppoe8eWxgdcxL8QP4lQhiowt4R1HQTpiZujEGYdvRxatAmsVfbzu0d2bLWlHjiw9yFfgY1XGP
GUrrGDb191XMAsq/BpmHTTDivSumx1Z2sC6TLICqyTMw65/aujywRtKbb78RvCQj6qnnASNPQ54e
Eve0hRV5UKXJGqCQZXujuWJFIOEMtks2NCJAPlfhjZWPNcjvJSyWB9DGFbL4Q7ncx9/oo/NdqRr0
4nIKqSXVyncg+V8+74h390dseoCR1MGyG/Y0qYLMH79iSQEgXo0k5l7josQfjIQcNWVWmlXVQDDx
wXtMWpikLQh9sF1PVlUdZ/UGgoOI6bsBOxfAShD3ZrE49XO09yzCJBsaqtlvpWichKL2n5ZxE7FY
UPk6AkJ24m1sXXsyz8nc+W15wSMVdx/j5AW7g2202pJGX+gjDAEnJPwO9SWQhnu6c0UYLbS+8Fce
W4oQ5+TfPU+oJcZuM1RZZu84Gt+F6z3luw02OyX60N4hsoidF8gzw0EAEokRNPj12Fsw2jPesDDG
6icFNubAlrz5a3euYrktZscesQLnPer9syxvLwZ4/BZ4fLtWKoHRO1LacPkD7+/c518aZlq4KxoQ
Jy9oNSKVnEDTmdbH0Z3MIUb0pdPqrT9dExk+ofepNOfgqVdY4sCY3MYhcYe2QMcNGEwuxmkcUMob
o6TvBT/6cwMYjkY5EqpjAfvQdr5GxP7+VHr+ePJIGcOVcHnHSCdujlwLexIoMoldtOrrcIchY6KE
2ps45DwjPXvsiy3jINssk+rk9O3z3y7YFLUvQShiVyvzepyjn4UpqR4pH/8nYEyU6NiunubYBLYJ
L7mlLgSfeYdWzwo0BhaY2bCuLJAnTwZ1VusI5as0LtlsLc6E6U4GoT/hQFzsIrPWxkWLzivDpUsc
HjLYxENw6cOjWC8b7YxRoUbyjvm7H0Jgs+dZhffmHKQuu884lXDWXL9dqN94ZWHF4VFPtZlSSsPt
GGDxfgPR7jDuHH/hdcAUp0nxDZBuXEwfOstYgUjLEn/16AqPkr54jbK0v0mRgBedraaB5eiyJsce
JBcnCrXfDQQQ1No6hafIgLtSFwKeq+WKOson6TFfgnrhxd24LQb+QWySiuI41c+6YfZrbldsVRsO
ULgc/lESohHgAwNoNttoCG9kdgf0tiY7pJOzuTfQBMZYMfHP+QOGzYy9R+lMA8uy8bRJFNUvXYxO
eEjvoj/1j2kdMSfFBl4djkVsg15WA7UJVYIjZHPROs4yGGs6ctkteswLU4q4+j8lwcDD891B+1EB
4l7dzF8GdDbj/i5pQE+FLRRoTT4CG//dZBpUlDO/hLDpqPOYNeO+P2eliIJGykWG/hWRvDTuvNYW
u+Z5M2Hgv2K6wpn7y7q+ebKQKJMjo951bb8CbYqPmWcUpT9vwvu7bFnzYJhblhg3g9oMhwsRuPAY
AIsK+vydrU9/1axKjw7rgpndt0EUcjESW+GQkxPK8GRXEhe3Xeo56KNyZTWyt4CgRW2+tZyF/KO3
yWacDIc3dvLTu6dsmSRb/jTTYZurY5ujM7K5ssbDZryUFLlOd7BM4TerIqEyfjU6GbWgfXLRQjqX
b5b6zNlXluugzobZ7MmA7oRyz8axD7AovKwwvU2gy4vX7wOeY/45SyEw/U832dbOZTtV5JzVQfzz
7WezbH9HNjMmegCLPrFnggzhZUvVDuUq2dOMbICk0174SS2EdUT9unV1pQ1/Y2omRq7GT9owd3YW
W+SrfhmVYl7Qe4cDU+U2l3vkPCTUftlWA0NH3lFG9xTw/VnsWVpxd5SPPkw7qvMMkdLgJr73By/b
C60fFoLTIXGm1k0Jyzovj/tlbu6J40Jy2SosY1YxAy9e7NYJS9xkM4RXPpZLBYINYoszvSsXiOlZ
IV+XHkTDcBFA5oArjHeAXa8mUmKvnDRxHhRcW6MdqkPYN6E7hJldpHKLq6PjjpZ5ZD5K8Q+nCMNw
lGv/NKlsPHT/HDRaLl1RlrBO6AfnEaDPHvNRZRKj4rQqrhqgYf1DXLjQLLht6s1WcmiC38dom7aI
f11uTzZPDSvWaB+kA+X6+6v3O5+3mAnu145sRRSpDGl3s2gVDmPpLafQHP65TvxTIj3v59w19VWm
J27hs6l80JCnuRsjJTxUrJYEKLbW2vnHV703G7H9bAGRql6GEFmJWdh6FuQRqgeq9whELDhIkyly
ifFjglAgUz9hc4QiNG9Z7a69TkRi+Uv7QPbMXdfu9JQmuK7WZp9my8D9cGj75R52ww8Bml9W4xEL
+9KHDbxw/LWDKULVsZ96KQkanINmFQdCYqXhnCsJZ73/P1WQbKrUR9PSsJZ7D/s/Qmx8bkaRWB7j
5D4q4PVYt8p7JgOx6XN4ag0laum34NvyG7rzTTpCDEh4UIvlvsnG3KctlFEKdAbehwI6D4GaNd/T
hDW58xdIMUmDG8Ws46Ee1Vp2e2vPx+5PXutYSzK4NkPrWHJy7poSgZMtoPdsemAqG4WBmSUJXmYJ
JD2+P3OdR8NnJwHbksvciTHrY2xqUf1weRlwQIFvKIYCrk53XHxiT0Spz1ppvd6uekm9tQRq2/7Z
qQNSxFztHHBQyd+D4QiD6fK0Tuh4U0k5TOUJiAtERQ/9kg2Eus2BG15lTcu079DxAV3sC6XTac1b
b6pKfD6E9df7SHtvMoDD52534HksfyY5x+GfU3RPVMocvwO7eDWWJDlp2BgzGjd9pz+MWkRsDIFO
KwYseDO1Sz6pcc1jhbgeXrovt+crVWabQklY0tKeuPVRwdrEuX8dkRCqfif2+c7sWKe578aaahKo
XKF4piwwUim0rAsk6mAAE0ZCz66TY6dYq0kJQrgcpAqs7Cx4SIDGkDqq3DYWqV/jZQgg+gBuVtfs
8BKZEtF2bz1kCHUe7vW2M7rAOQha1qRXn7hxeNUNSLTDijGNsgNDvyZOKPIUlUJoyitQm4m/rDew
rigwsTMTQjgfiz0j2GuUb+gP4JmQ2Uq4GYIvGKRxLcsfxwfZ9fgUHbZWFqAvT23a+NkrW5kYc1HQ
OsHz+TVY5GGQqWJ+X7tSaOVCJcxPEUGPdUxIgnQ49eWYef87xfucuryOQx8lA4TvXQJExJ0F5V0p
PXmNi1c8Za3yATskZCQXlS+DDwb9ovStc/OLHYFB7vn27kD2TAsvKBi71k/7TFr6z7nNSckt6Ush
NKkDAbGAkU37K+Xw/ETuHoONSI0tYNgw08+ec0zvx8JMUPhKaMYop7HvSRQd8hw5mToZnsztrCA6
Xba2hMFqjCUbcS0dGKYWdEmieP1Jzitj5jxM2BW0JNqViDfjfHnIDy9VAU6moLXHaUd4Vjqee4oU
0nnFM0LDuNPWnHaBzRa352xLhfC/0NNDsMtMrdx09dMgeIXjEM+TVTvDg+jqyE1AWZAYA7mHg25m
iUdMTvU6p+O9vViMdmWChQNfG6WMkkyrTbPUCD6IsGAwlifYzlRyEkzbYyLz19Ho0j7AOzEsZgmW
hdbuPCEvdgEhaWFxJvzLIqqTP7Kjmjr/uM0TY+PneNHeM7UDphqv3JhW2wbCQbtwaE8IcFsI5Dyc
WDJ1BaJ2SsAvJHqiPJmCOxrnIwkMlHp1i4bMcex2Tq408WB0Kz5HVfggalcdL2WPWtpje38EX+FI
GP4vtv0wkQftDD3bfQwZDCrvJOcK79FuXiHclxI8VS3Df3WJN5kuMqIvbn0GFM5rF+G0gYNmgGoL
SAc6xomdGahHpIGhF3tz2pU0alVbPsSB0Myc36/fkSMrttOGSoNJF2HH4ehPoGQyARTwqPqbHSLu
F4cDiiJkkOnzBkmzElPMMTxJ4I3QjX58hw2TPYwSLaFCHbn6t1FiZxiDNAlgRHxubYwLh/eDA8Vu
mzN4JtxrmNj+pMXbYUSjs72lRKXwtl85zJB0Q5fr7xOy94t7CsSkK1kTKimdGX3tuw+rgbjbxMFl
wbEfIRrGt8d4xzKaEXxE2gWPy5VjSCXJxdPTbx6MYI0+uptn9XJksjKBHMQFGY5WJ4zJiEE4X9xl
tvb4bgxtJsVhDeNGpU1jHGOKEE58UOXU55+uS5xFvSfT+fn6AMIfckWfT4/mjHK+h6tff0RLzjTl
tcXnaD+YlqCl4oZhTHgYo+vhrKbYb1/F8G5LTSMNHCFlnoHZG9peUrScqWzZ2tWK4TuHeQuQhTk+
8FoMrrnREiR0zum7dNXxJPvn4rl2c1IvZdVvYPrpBviDk2i/oSaIGcH2bGNxmRO5MGo/KJeEpDxq
UZ8aIxIg7fTDkV11iGK6iM0khuaDdDGRo4/thpM62a9F2h6F/3BA00XUyf+ex7YZ+RdQuqQvtfH3
MD8O7PbHTqaXLLvIbhHSOZjLn9X3cD6OJ0nvoI4UrmcqwtY7IJ3/fYaGM2srRlpFLGP3E+rMuHHW
xokzBeNsy3MEcz1cMu5txoCvKMMg7XsQE91CLa17CbGkVkw1mpFqNe/pH0Q9IdA/C7FsNf970jOp
pnnl+hz3QJ7urvt8qPuJvd+DDfq1PP4+555KADwwKCGIPzEOKzQT1vdkSrU8QckoeWyy/6O0Ya8W
YQAc4GM/P3rPW8/CLwcbEJQirDOH8OQwLg0iO0dA+r/vRPrDqyuwWGRfJBfdrO/R7qP/ozubNw7a
B6XyuqcGBS7df+eyq4v1nQAIuTgcPPiNBk/ZpLQu7ueK8fT6QUHUUh2rciymqZ0J0skVHJyOsx/E
ST8UU/vOVcT6UFv8Xc8C1PyCxUyxLiMEXGu90dUvUhxXSjb6so2Zz8//EbFkKH933My2Lfz4PJCE
tTwZGU/n5uAOjik8b0CnheZ6E8xPXJCXXxBEnA9iuSeaein2VfvOBWn0WxJ0C9jWt2L7E1LNUfpI
xkQ7MQroSjgUCqPqgUhQ8zx+jwrWuX1ReTND5QGdpX74Z9H40LI4ntytoae/jra3PAeoToLJlBjd
D6pKtd5ucrvdJbPp8dcOojKI8ta16eIxAc2UXxbEUGpbUJ5HxlhpVaAeRwn8YKB+AcWFrF/Q3r4d
Hj4OMaMltYCyw7NWULI/iKN1Rzp+K/9fqq40ihD+TLpKysUFFwcHhthFCH7zqXuZ5NFHh16Gn1Lz
vpq0tsJIcH3SQyRADK7jOpwvGW7qD9vbG2jOq8k/aR34sC3O7aE24luUPgjc/Yfazxf+Rm3FAXxf
9XK8Gj7GMzHmWma10dlj+F/YOggpPhNC2FcZ8UIMEUNch1GE4qEKkf8KX4XkG8zuth2kBr9tIUKh
jrmNRBTJoyRHwwb8H0xdSnYPjv0aZvmwZUdSK4xXkT08q6ndgOyQUI8PnDE9LNxila87QNYhQn/4
bgn58pGb4NMMbiCh78epWMTKoOIbTbFw4lhGCaZpjNwmXpigv9Hm6tWvgXokcKu5fAW1+V1dA20D
8ahtsIezKtFqZvx82dw8tc3Flw4RexHQC8Dhl2dAA9H1wpRIOCDj8scKLpoQHfTO/huZj3nRvpmf
NFPR1YRrcrq0AFrvDZPHw1wMQRAwfvPf50CW31MjsmLhJfaUhq4vlxbUdYh1PKohNpSBJjE2QE5G
eAaAwcvy1NAHX91UaP+wWvSNWCt2yC3Ql1p7dCMXGa02rZZzsGTpXGV0kYePB2hnGlZsyFwPcqpY
IlN9JSDZc4oc1CltKP2RPlxPzRM4I8QidGZeGTzwDBR/xXmL5uVJm8EBR8/rNIzoKunBdN1b8FXZ
P0WZGh1MYMXSGVJAsJL5uDIIVD1ZJOqSuYnim4pFn9R5WkAbxE3Da68jdfnta7Comjb/X3ubBa64
iXJZm+0A41yP/dsSX2EMIEeNrlD1+I/xjJSS+OwdMxmX7z8IBOVpwPSMAmfF3wyfOpVsf87MK9H6
pmhJnhUWXNndjr/DjyjBLY1xDaFlxjjQUGFwkstG1mmk4s/XZjxM91nojIoV1u6Y9OqRB2V8RbPU
eTAsFclCPbHutfHS4oi5tFp6xbW+aQvHXv2GhJ+SQMy6tCDWGtim3SDVTybP06LkWe7VOtx2SUZr
1ntlx4+66LEB1cfJSY5yMI6KYJvDxGw5WHROytwN8lPaa953RR5wgzf31BRs+MzO7jy/lA2MqFdI
lVbj5lex9XfdfQHsCRxB9UmPEw56Za9WWNdL7cICJWYWHAmCRDXQgB+hvFten5c9qmyEBuHwOpmB
hyJ9zTeg8dvTrJDIulo7dD0IzXMKxBxs6OM1ToWWzqpTGops0KhZeJvEzziy5yl/I8wEYWbIW0z0
wBSEqcnRq7dmw4ophtmXpQnuB697hev5QjEbc1w2+Gr6ckwH19aOcLFoOZidEg/2rLFcj5fpQj4m
FAYI7WGWsIlKtEQLyDJcBWjjTa081RkRtcRojjeJKoRKQtNBBjj5sCNqokgd/twII1++DVDiqD1D
hIoSY4nexMJ+J+yjbL1IfaXZEUYq1Yw1LVtB1Q7aRp/g8d+sDf+fgnhKv+0HduwMFZ5MmAySdhaY
Ccf5ZyjQ1XJk9QNr5l14y6NuJIsqxa1Ye4xlnVpr2cfMTA4ufBtrrwqmZwIrBvg1xDHuF0vIl6af
qlG/gi+mcn2vKdaHfCWUXum9on1R7eicNHmjJB99GJLPv2oCtDSG17bBylseBtqO1lTMsRi3/aZZ
5C/dY6962LR3od3IoAsfY4KEkpf2D+onm/K31WTlQc7rW9nnsWDCUAPf/AF04nR12zqtFZ8pQxKW
En6hXO1EfaYdHktiqnXJZ/Eliqj4dtii3TNzKDqgTeiwVl+Yavjlp6dxW9hOGrQl7ANEYsXDE+G1
lWxydqvy3si9YyFj+MyzmcyYsdmrbDUb+LfsMcQGzeJuSOv3SJP07PIjeNHtV2mQuwrW9LQa7lSR
L2T+HkkdyhDIFs+jhhzS5I8ku8N4dOb0mE7/nH4MMGn2hfaWjoPkTDMtig/uhmHU48OJROR+hytC
bNz7C367SPGngKYYRFR3L9AlpHA5aiarEBQiD+MMApVpj1RuXL7KnX0Q/9FhIsfl+9lNS/ASN/T4
E1F3MrPAoetY9rWBAJLrtJhsMQf4/u3KJ81PE42QtyTj5lpxrJ4nvNWGXasvpJSF0JzTA/wLsGbD
IkzyeltAv20M64lMCBF26Pkb0Bc0itYrdMsYg3ElmYWjDu+cREERu2zUpuwBSvJiGi+ro56HDwOZ
7P0iWOnkCHhH1xW4xtmfQ0hQVgcsmAjUUlin8tb/7TCeWDYciForV/lvLZwzlx2Pspmm1nMJoXPI
d3BYPKavohC/IBsF/3u/6gw5FC1rJbEVlzIzlLhNYA9CcLb4GPyPwlkTIv4RecBbgh4tPifFZbLE
Q37BgU6JGHWk15Gjai+ajbE8Jgei6JgSM0occe/dDTZ+b/j5TnBPLaN2a1YmyUbqJ5t7gS0z9wcl
n0m8c1NI1jEF2DHYocAUdRwQFqZuvPHUQoQFsgh1zBfAzOXcQ2tC9ht4yqsShJgLUrMlor9l8JM9
Nvb52qMsaZII+8veqE8oFQKspElbj1GW4ckzvHCGNUMuP02YIxMoo/ZHqGZprnh4EhyL6zEeo817
c6T6szW9GLNcBRMuy4t7lFG3lJ7i6BiVmlg14vmm2T6NeaRhKbdHV70Vae7Bhb3pdu6U6ZJ3VMJs
/02tJud4Jl6iTrCyF8EdrFs6kFkFaLJSDdTyfNvDxB1HCBqtbEWee9rjj5rmE5AJmXInjDZYUGQA
jvgggH0FiVgPQsfn6hYyVwaiATg0oEG6pwIHmiyLh/W49L9aGqkotAQdhJNVfC56uzs2QxKX8T9G
UTQPL/Kvmm8JRxa6cvCWoTW5C4YCTWs31oq3Fkv3nxh9FdnDP0QB4F7MPTrYOsn5jLiPfraAQNA/
yPrEexRlFxsCDR2Y8owfLOYkakahV2c0x/v2Ngds5sH9eOK4ziT7ZFLafJbMb/btqeRruRmJ8YLA
KrIoGqTF5j1ojLPje2xbqDq1m/ssy7Tmjr2Sv44NqbNjVeCoG2C7KuY7GITrvB7XWII7XBfxc4Ba
XKu8kDTesNM8yUQThKSymwZeWwqNrEvTa1owfzY/QVSepftNdwH54qVMy5TGNq/RM5OxSDrHbVn9
KI6S4xX6VSro9Nn3XtcEnKKq4NrLIfhXWHo2UgJ9kO4O9EP8Xcjh7yzBmjIrf3A93P5BQ1P3Txhu
0neXnblrmQG40y/SAXEkPGlkKySepPr8LxmBm9/X3UWUZ0VTu/pfSzd1B8VseV1Q9PDP+OYiiinm
zA1g3St+1U6ITTZq8EazYw9bV68P8+0udRVQJdHu2P5chWK1A9fY6IOn8QvTwm/yQFr/FlY+AHvY
vP027CiHOnMRW2X+Yjy93E//zJNLHZCHfS/0szL2vYd66HxMlpEZeRB8wuU37Mj/qGDTy/PFQFKJ
gSk3Cik3SWYHKcqWb0dQde+NjXYDRoEke73U0vAN5gjPKS+X2BX63iBXdiNlnz9cyH1CBSZR/Ua2
uqUxaFcKoFYlqpiwfDQdRFTfAoo/wcquDYPvhkcTBLUDZaH33EInprGUkGnKYFTK55nhtfGDvuvo
WysddPejQTm1rvDGtgwHHyEjpGOJxB1Ef2qhTgcBIHvlblzTRkzs8bIEyN1qu6LHH5dVlInoQIcS
cHCuBJv+5ti6f44/aKPw+9JwfxpZoptSygZX64IOKnPjo2R6yuod7D2nKRGF0kFP/KwQnB2QjwRN
DnCg6k98ZbZolEbv8q2eP1BqxvG81vfnDarZiS4IgcImOXFcjTmjlj4nBaGkpKc3tftdvmXoxsMs
hGszFmAe8LsDeRa6qyDDiy5FIftWMHntaMYyMY+Sn8JXCaGlgVt1uT+ulnzGhjAZeIX7yre/CBzb
RcvLpo0uLDawLVxWgS14lHzt9nbaBn1p+Uj4tbS87Uhw6cTKXTTv+2gpF/ggM6/Km0JfGJDSGH7/
7+9w7Usa4aR2CmT+r8ZoZM2uLUg0k8HrP+2W8JE0J/7pw04g4JY2td3nUyKxOoKFNJltrJ6ujXV7
17vYZQ8JmKq+PgteFBW/+ustaHkA7e9qNovByqiUHCu71ZmSgDNNCYKK/K7jqdaQP3Ay0PO701bW
GNY6F1WTjYgUj4MZDjae9MsWTxb7QByZlSXIztFVwOUOwjuAUvVIsSpDKBTgUE/tpth9r9kB5Si1
QvpcbmkoNRXJ4Mjc7er46aWKj8bVOYwHqF7iQ+eIqaPPz3nwTRBAMd36vctykDILClY88v+r7YDB
ZdBaJURgtD00/fWlxlU9YdlTaltO5ylqJDxQsml1bpjO/Rskz5HnUF++i7+6xtXy1jx3o6WKPnFc
2y8BDfCItio9/uzmmAUvwGi8OTN/YbaIFZcn9NFU+fXzpGQyQQfiuJNdjTTAA57twb4ePX+kQ8Pb
JfTzPDZ1qXLhc/2312miZ1rOa2gDOBkxLEkk8R6t+8KDR1s/YRhXrODMzzb40CS9mrzlYsc/H/Ti
w6hvJiO8vFN2FVa4/yd5zWmewAjb5FzCvYl5tyRduUk07JIXQuWhDGHOXhaYNDoDuQTjdhKgiIjV
1WWqz8jaeCRQAO2vHNWKFR9z3gaDr3UJrvhFYQ1i0XQX+1PqazIzQlWzwecivRiVB0CTgUzNWXY9
zxyus+H1n/7VqOB4IJmhk/RwxlPZPqDh10GCLLGKwBwzadMcKA/jTM+ya+mNBdHAuluUwVDF6BaO
rRY9wRX8dFebPXeAJhd3TSQKTzxMxbozIzwNIPi37jdYSucTQChpDGtS8I4j/eWB8rWCkg5SalCR
hx3CctxqEYWzgaMSUUwjFeto1n2tmEtt+oknoIG4bIzmRdYMJioryvLhRQl2xYTIIl5GxyoyLTX9
0pRDBHJJxylogeDuqm2SLdphZ9yq91vPfoyWJRUngYYzNjRUgUxDlpzZgIy7r5R/P2q1auMkPrvC
+hwitmkGTT5o1ehtibumWq1rZLt+lxYRRyAUuPw93Cv1303oZvOS6fMhvl3rj8wVmoakgjD3Wctp
WgrfzqD+WrQo/mAQ/3803tBwbm/A4VH4h268YWU2AneFp9jR9i6A50EmqXenitR7x6XxNSZA0djj
+gX7fE6bAklNdXQ546Xy8iJRpmYpMDou8cqDmwe+Bm+YaeCYTCSQ8TM2udJh0y9V6ug7BkfVxSzN
UoDo154Qrhd06kphG/hta1Ee75VDwzBvgcxWm+JHllSVusqTk2jyetMa1zEn4CITISHQBBiqQ5jN
VKMrd3WbMZR+UvcBGeX83bOCSARFC8R7kdr7GEWN+JBoG0P3uiYE2+9j1wbbGa0zDp1C0NKUE+z4
BcrP0jrnB+fSdU1/GPWumBcnJdQpoccAaWyxSPPwg/mtQu2rDf83GXY/manlASf/E0wRS7IIVrPW
7l2Tg2ObLkltgu2ZPeuXnVEwPpFhcF+rftUmLu/qh7ueRV+JyY9uN3cLeKJcmESpz+TbyTBAkIpM
OB6UQRk2nDlhWzxN3WLYpmhVkUB40NTMUZd8pDrWtYikULekS4XWVMEdvfGTxnDcQesCVDvcK9U9
v0k3ve80GcBf/Fe++JSXlDYGNDUWL4+CYfE1o/WXkI2blt4aFcPvdNtGnzmXJJrOiJCvmOfQzBd8
RPHd25MVfP3HFa4UPqRpcknwAOIdCXr21vxLFCZf1BmEATMmFd6oJgNiiSPuSbYSuNRqOm6hcpwc
Tka4Z2PIE1/yl8oU3YoDdOTMSX82NEyE8pKMz9A7ZbfWUVJl5xepR7yp716dC70L7V3HJ0Y2pEAY
WSASBDluwpOh+QhcGwFqjETBgmeEvxaZsPyMc801GCI4iR8AMoPZoG5UGJUJG2vfLrb8U5gjPRk4
eYBjYGMP/U+kXT7+mC2AlQwPpKZglc+1AveNfJzF+OqMOfxoXfBxM4mqAWuit3ftPASo0PyWp8KF
C2byk68o2/eYv7ei0it3OjmaKiqUbSiqGlL8Cs55GASWoxs9KEJcNRSGeipCDKo067jEOOmVYNfV
ZiIpSLvJJ7W3ZSKN/z35U8pLbN52FcGyYekOw1s1/UIP8wwngFNK+ykEl9jc177/LpzdbgXdD6zr
NVsAf3BlyMgLvF68S5h/QO5BkrTo3ZCPu1z961A5MwN80fZ0IgxLMPnw4jWuBC2CsGf7FgjR/1hK
RSwDL7SiD6MB4m3iB9OxSEwofEwLjrgWJax+TZDYToBSiRV4aN2J43fAXWe3jqbcM5LITMoP2FVf
X0fDSeZ8YtpVL6SQGp0vzW/Uqg6X8VSFbnvwwQVy//s0AkxYdr28UchuXiGuEfdCjqKWoQ1EZ1y1
WvngwW6BpFX7xLT6X4pROzzcVejkIGECXiMrKNoF/OkjGwDx0MTGHrKnMcrqcrdqUMPSc7eLApyE
sQWdLPU7wxvsLSHZ/iHLrivBqm7gW6pBy1Q1XsJDpHYtdYH8FdZDa/SKwe6umkvw2/riid9YaIYk
HjaShMofYQEcPIizYBGiNaWzSqViqdoQ+psvgePPTpuiCa7sB6gSKUx5kNrzuoLatJdLgJTQapDJ
GEUlj83PRvTt5jIr1b2e5T25jBQ/27fKhDiMgaEDtZLFZIR9hEvXkaGh8dGNraCqcIeh/PXn9nS0
HzwLBItqdb+JtnTPmGaO/qKaRb2hFu/5B8RxITwlqLf/w/Vt+hLLS2/lLUGaBqLv5jJPCWhaElyP
aN2NOelNJskdcSEu49OMzF8dJySos1WSvlaH9NFAKb+fDI/JI6PitZsy4d3YEWrElctkzITCjiSC
QKx8uDoRa8RmOzX7GdJx6enlHQzmURLLtrV6C4UPfBEedfoqK7cEtiWBByH6gIgiza1EQXHzPaq5
+vzgdMILnhMT/o/zqiPRjpEBG5RZa8HmEnc2dfRi5XdC/xSzkcV17KJg/dc0urwcUtb/R/lZpN/D
C0j19JcBwLiUM9HJKiYMVzgwhpwgKgHoKMY6Hl05M3VGgju+llLTcQ229ARFUCqfi1npVoOw8YgR
gsbiqlSs4HfGJsenMmSRc8Q9wSfujAELb1fJJ7ciPR1fo+m7DpxOrTq/l45EaaffpDxvyKUy5ywJ
SY7serhEMdZsSio8mlsJL3URtLuSqZGDUR3MtGTvWBcTNbgRXL6Kb+I2B+AA0F/bqC12fYgsxQwq
ywGz3C991+Krf2j2U/65lnzitb5q1lfu3EEa64zvet2g0zVLm6TlOPQbarwvjKDuJdJTUdJoIVol
f1u5N352BaFBtif58r23Tz0FCQ3M+INUCKUvGE3YPpWfuiFuPG/QG9Kbj1e23dGOOi98pfW9EdIV
grGEZwUMPoqGHtUeDO+vXb2GKmk1cdNw1Gqp/erfXrvpK3B5eqWnUwux6bMltg4iqdiRLUWDzv5y
HiHP1D/iWaYKbAlJqyykDdj2ya2ia9KDaS8sfr13JXTlSrUUUp+rQllG+dk2QoNea9aM4VuMKjU2
hP0tjDwAlh3X/yMgExa0lRKaRlpiYqDVR2ASq3mR5kqvac6xgsX4W7zge3i3f31COAOxzDzSClFL
6hVV0n4L63hePr9tZMEsFTDpaUBKGRonvzKfPnh7tky7hzSmY8AGjgRorgI9aZlP9wPQyXsLPmId
Vk8pco/A01msws7MHrM3xI71+kQL1k1c6jDtaGOE4PTl8XadTNszGpHH4eZtBI/3aEX78gOObxrk
KmchTI6z0cYmMP6krvEqfH8kb+/sxzrCDpmfqZvSF7xIIuJsKgejcVo4IbJS5wK4aLe5L04S60Zl
Y8UG3bjEGWGXGcSsuLtrkRwWZtTjn91ivVGSI5E5GRRerb07xdI8DDy70Mnszr/JvB4vazgGkiB5
UgLeyZCeY6GuNciEit0s0zOX+trkAQEqLG2lk1+HmV1ukQ18m0LfQ4aPOyUMW4m5/cFEEkeWH2wj
Lo7KMEp/dlnlsms08SLUs3V+MG6LjG8ddXU5a1o3ELmaT41UYEfGhvBLjq3dqOu4Wb3wUpdmjooc
M23rTA+PLb7bOR/k25ET6+EXd++iWUjU1lXzYq4XbPQpy2lDAqGnqIxPlPk/tpJWu05szJS2zGx/
XEU6SnHq3gSApVhaScES6Or6ZCo5FeOWc0sqK7mK+IzQG23Dbvexa2+D3mjIiR7go7O7qjpRgNgY
MT/d2Qk4bH00DhPDSBaGz/p5epFPqpsb9vf0rmaz9XcFnLYo97uA65uMUaV3c1zM2NmTnOz8WkBB
TITap9MxO5raOnU4NEh/GQv+dZn4RE4Q7Mumn8nGcjZO9eVV4aPJXcCM6bXmK8w/Ha8UktxSE73v
DurPcGoAOJU6/l3c+67+ozJfYTaugSl8SZMP2x/rSKqGO0xAMe4pNa4c8CEubV3+9dDiUhAVHuCS
QXzUyH68yz+TaUczb8PzQQYDrEjQ3q0Ujk01HRa4qlLyOqFwq69Y3FeszNpCtqdVI3H9W6rE4vlp
n2f0WmfwS0d0l/zAQpeKzZ5ezsghdlTxd1ZycnJ1JVg8QhmV1pCoAp9lpDAgxp2UDq5y+HFp5+dd
HAWcAbWqhql+8KP2eBUIEiHmceI/TE00bRmensiy/44nToZNlMTkPIEvV2ei6gid2QW+tvf0U3iJ
SIeSmAe9SeVDoyDBu/QDL31KiJ0ARYd/Tb06f9/h+Qzvr7jHbu0g955EP181acmESV0FQxIEC19o
BTlq8aVlBpeo8j8V+P4urOhazxtkjB7miF5YbjCMrjfGJlADf2Haw3r23xXnYbZhZMP11VM1gdYT
6y3qYx/votfN5ycz90TfVFDm3nZoNdyZw1LoKsmca/DNEsRy6UhngKfvPZAVAt7/0/T4tViO/IOj
hJT3ZCOtAR8qP2pu13HvR5CRXfcVMq53yl49gGWNUJjBz7w+1JGRnAHN3xxth22K17cMDsrHDOhs
aXn9HooDbuVbzewyfmLq1sN/a7mrg2m0/WZKpTcb/5ieBe1QkiOZmuIvXnJzLfVcUnKNIBTcMUp9
3EvbTKClGvR49vNielT0ZF8VNDQCQGBsILy5/0dNZfJX0gYYvcuNoD/yGjeUB4vFu8JBV0URWec1
49ljqIwQtWn5qGOijizwN4wIjzwni5JC0mcR4GafQyDDSOO66g+w+weWh7O4im3USlA2BD4Sr/6A
LCqtdQPlK9+kfR9F3enVGA54CKkihL0WZFjpNflbjttOmp1w/eBciwldBWS54rqOMki4MCWRlrYL
CtoAgHuoQXAeA9tmtA/D3Qmjk3FicMrhIjVk6mDv4wFO0SVYZLxhtNhKEoKEWholg7tSbXi0ET7m
KGaB60lA/63U/w2V+qj9IviBE4xir6+H/y+LDY2WeBVplBtAAqig/ql0eYI/4CIAWxoewxHbbSSj
380+RYUBOw0BRu5SHcEUfu5EmPIS4BknIX2/Y8pwe665mPfT2hRrtPm7YAyCYMusMsyYsF0Ifnpp
Q3q6gWk0tOWYIuEEcbiCJFDc5beuPjFrcfazYI20b1sraH3OcWN/zspqxdhBKOeSgEyCrejmGj64
czfEkhRKMb4ef9+NSr3lmlkAh6uaR+Qh/E/8K3kTgK8lGjOed66AGuaCbLenJrBkUK6vxfVxJBvb
57KARZ1Vt8HrAbzBB3NkwLWNn9YIoMRSjWQrla6bc4wC6K0JlqF14/KHXKHwY/kEP9iWjK3GgY9X
BcR7UuZ31Ca+Oew98Qk3ZszEjrcbreMGUYfHZqSEx3IcogAtXtksxiBHEt+aIVM08iVlDQhPOdgj
c89ch8xuD/r5v2G3GfB00PgwVrGwUO8GqZ5gwqYsFMXFtVwXvRQqyBmuhYOrQoGe4FBtxyKUnHfz
6ONg7C/jHkR45qqiudP+TZzS1IF58gcOJsIxwYWAHfaAkXFBQks0SqwxMXjiOr+qX2T0hYYAN8kF
wpQv0vB+y/b7DZOVVeo9uEP0x081q0099YC/2bqEv3ZqEGVPFmlWYBw3gsxyKOBIloljxoYN/8zc
yLcPzIbW8XJV2pKMaBhtEoOne5aOVRUko79z0UDPZSMlyAL1NvfD/GWn/nIOIoY0zCOYcOiWrSRC
8he02hirQD8pc/exSTZW3F/rXo3Ac/L2U6rs1ezJmEZupljR3FMF5Ui5ebXHn8kv4ETJXBp/kw7C
o9ZWxEQlTngPeUUata+gPl/16N9U6whe9SwAzOiCagP6iDHtVM+loNzWqblI4IqXEl0OICpT6j8y
7lc0XgqKiLaJXvwqxF5xD9jxkpBHPAeqwc7jRdIpXb9jfaJLTsY6w+YSHfgEDjh3L3rjbxxGqt6K
lcOZ45BQE5NQEsJxmzfQeNz2BwM33LuKJnWchhWFMUxvMSDauvuhBwVaGAxoQGBrUh0r3/jq7jwT
28FFwf0FOZjXnjrb3M1VLBQqwec70sZy0EYsP6dUvcOaE5SD26JR0kHpgeF1gjmznY2VvpDeVhZY
GHAePTCh11W/B77dtT6u28GJdZmQH6na0VD8Oh9vgtlXHGUc02e4hSF92cgtZ/xXbVVe6PkZ/DCJ
wKpRI5D63g/TY+klohVAJ2r51g7KvVRAMJMXX5aXAd0rLxpDHtNIUaMYbnaGk+s+znU7jcqBtB5C
4CALQyJszkSioLWMcA+neIMy4AelG8E1nUwv+HEJ2c/DXt8pB0G8t7pv/OOMrOgI1k87DkwL4C/E
pxUvgrnp+ffO3sGNyGBSFkKKiAllNS9cMENz6p/le0Y1vdfNDYyiIca3hwQpQV5t+A+Echz5XH7H
HBoEIf/66BnmLqr5jQulYiFD1WoIoEnG98GnHf8GgHQokPOaxUVcobIHWdgZzaopNWqfMMLZB8V0
NPLanoAEopQttq5EoslRCtjAPGmBrgytcSUjPgIBUlCtvZ/ljXOIp9K6pZzGM1GrNJowFmga6iUn
wdlohCHUX6ggqetj1ET5FHp3cPpOIFjmReCXZQXf53pZlAtn1/M1gA9HqDeRF/G5v6EFww57mxsz
O2KBZTUAYwdnoWCCuhGt8V81q7IJE80l3i79GAqBrjBkstAMFklRZI5FLHdJZXawyJveYlo6gD2i
f3ttRkB93v92GfYiuS/bNRbKSjwiedowdNOqW9T5yniNbZdlHLencWmyWshS17mw+KKpUV4KdyMN
Kn3cPGTMbjCbBP0sCpGWC4/Gei6krY/uu8UYkW52m1dcYQjBq5SG30eTvsGM9dBlz/4Bviii4Sqo
gTiqtNfBgHyynMjBcMW7Evf8RUfQBoaN5iva6FyEPwZ1EwBIP5YzNNX+t/GyzcCAiJNSIadJQ1ha
E3/HRCZYqQCKnVoSJyDuTk5swDGQzNkDv04BbjIaHBh5XhMjtr82KGLyGyDjosuiK7jRHV1fbjqQ
J0ency7e5iJaOX8D1uKp9x6Ej+4qa/8QBF6fSWnnZ4ad0jnsJ/G0EzD9bugAg7HHA4OEF6E5VGNm
TBThAOuMdbeD2EqMf1fcgbLdd5OM7Ol9lYUCAII4f6fNxg83k7CzxClL+vFZQfLYoUJbq86xsBUK
K1jojia/+9sfIFqEuvs/D1IrH1V6Z1jcG/xEfKhL14FMUhlZdeDc71IUBuXrfaEDLOY2MHmgj0cd
lIL0mcd3C7zFDCAY3Vl4VSHJcnkJkvGVts/qZiRE3jr7iZSumgjUHzL4jPOVVnT3dqfrE4Cbb5n8
ptD/jeR1LTIMnBc98lBEnvr4EulS0hC4O7QeTY3iNbW+tRRu6mu1yxgV6HiGBi+Ncw5/vD6kJ8Dx
5HLtxovEv0vBC1iZzk6inbVHhaMjY2m2Rzjt6LhmHDsgrTCS2Bp2RtbfsYXUqEh+QyXoXY7bTHgI
e8ZrSoAz0xjfZ4LGsx6mCTOh3keO7lBLFRXRBt+9s+/t0Y+zce/1nvqeBFExm9NGN2e39m4OMDB9
jDce8h3iFC/+mEIX2du07wzZfS3FlIyfw2zCDCfMzf1wTLK2Xxq5yUwQwqOW8XuSe9Z244kzsgeH
M7G48LeX8Wv0mZBbaoJAJ7faihf0o/58a/UaRTwD8ZHnzUV6UPzQn4HAi1uJag8Q6HYZggM4A3Iu
uqkp57/3Ffd+2OfCiUWmXLur9+njbuEq4Ks38LBUtxousC2hHe7JQCwMwxXrbtsBKZ+5w1kFgOwl
aCKVCIOTs1ZX/jXyqCaC1p0gFjFHppyFfBxFIF1Ri5Y9x6Xyhc9wfULzBXbhYrUcrRFU0GN7vjir
2hhr0Yvlobhtro9ECsddY3PN/XZA8vC6wJ1eoPNKsRPo2rpE66rgLvAAoUMLn+i8cQN6gqoSkomw
gloTfyc4i6QaVtmwbfkXNls9oauEzAF1d48/ThQnNdxGXAQ2jTnj7fVN6QqbMK8ukGNnfDkZr2Pb
jjVKaTz0krkMcNrI5bUBqWHJbfseqmABx8eFOCZKJQYtdM2pv1D3AhLs7o/AOH5k1UotOyvApfEP
JiHiCvf3dr7I++LpHr87Akw/wYdVpOVynunDE2J7ieO0I0YjDRDrldkR0JoN/d47g5x7pM6mDBH8
/+kz1tLmcdjiYS8GODd37j4JfUsAL/NPCNMC9CYlqAVXTtb/RYaSfELyzR0ot7aXxj3ivZ3Q8kNj
gM/F+n7Ou3QOsUW1u9SUmNN/68qAgkPEHrUzvvibVHZ5FfCXA20Xd15GPcc6sQ5kGsJqx5NGAkrc
SwJznQu+Ar4mES3+hhrpDwhtgczLunEZ3J2eiO7wciBaHZMYosXyShcnhNAn5rw/t7nKMKUI3eZh
i7S8oIkmWBoJ9IaAaiqGqw6S0oYG/GtJi6uy+wUdbITeIM9Efhtbc2YBn1NqmwTNHEOQuM0nm6/V
ADSGN8LP9HjeUbdQwmyi2Z+KZrsLbUXe+5G8ExJkMQAL+c32gBhI/CR+mM2VcZu8YCj14otRBneE
d0aN+nu2KMb+lWLeLN4UofOYPLSB7UjmYNzIItzCl/lF0EwOuKMrrjvJlXJrm0HAUqD5LlEKx0td
aW/Nz1BCIXA45qrytnGYHliW4uXV60NaMgQ5oNPOYWrL6miKtm4yONTSZArrbNYNt5f9yf/gMvD2
Ar6qZhc5l0dmd4KG2CVj+yk6jYLwzZppohTKe06Pp0hSGNqfI/EvICMGnAHjghqFq+LIMl4OOUe4
UfI6eCzOsavmBW9UG9WffLNWHtroTTE0FzheYAmO8SNGEho1jQFy0Jok/Npgm1P6Lq1LiK1mneOO
3EDhK+PU9jTz/PplrKVZAoFY/qzvY83qDene7XFSkjecJ5ObuASH3oqBvm9+/su+UfKrgFrxKpi1
jbiUMA5SzNWu1JX/Fm0Jj/GO9Q9jm1fdupbfxjIGT4SxcoXBfYBPQtepu3rcG7nWAS2g7PRY6pcA
JTII658bV5btnRAHUYV+ouBsH/9cKILqMteqrbEp/XKPZMfY8fNnEM2q0VBJ1/6fjIEjnaVDbh5K
Eux6BsQUiQ1ITUVTaFez0H+JuP19emYjrPLjRiQDYKbiWr9WXd8i8YOQoqnZB7BShLvG7Wdjq1CJ
EGubSwcEDWNUngOtVe8YYO8bKzOUy6XBgwU/SASnxkk5JgojhOScfb/p2i2v8of7pG24iJZMExlD
Ocu3GS+PQdpy6jYWUvovvnMfPrpXHo2nEB8zfc/d7DW4rAqpOzCcCroujIJqVWD1cR5CHETUeRfA
I0sur7LjmfwEZ+E4nSDUz37n9tqZsITrolFz3O4ktd6akBGMU88+/wMuRguT5wyIiYpB9nI4YDYl
S6MhHQWg8HY+YZVU0iDwusEUxfwI7a78UsbGFv/0mFPKwhzi8kRZ0oyty1FpgnheLl9zbwZ1aXME
aM2s/3O4SG0ekXlDiMw68VCu9O6Fs8nOjdCLapXyiJuc3SBtyTW+htwIhAH3lMlkBz5zJOSaKLxh
IfvlN/fhte5j9sG0qmFMXBARSIrzBEWeXzcvmVjVpVGpyKfGUpYgFzpXqfgrvFXcWHK24A7l2B5v
K7xH8TnzezJ+Njj7rt+wWjDN1ZpCOZaUJF1tzCwpWdPTi9vBTBjFd8MMtdQNoEzdn3M2rHY6e8Ux
MB90XSZ4csn2kfOCqnLTLI9/rBYOtiCjX76sRLrkfgxi9AIlltWixY8aZ1l5j+eZ0CVUO2dI7Pbu
KT0FO+cE0uo/tEw238W50KS7HzzKCewWBRxm6FLow+fl30CsIhAXSc9o+Za7V79nPgwF5W/wnWP/
UYndhK48j8HGH94ENhTVTQA1Vzyv3KwGbmhWI/7BsTzEHvv+1aR+z4VabtF4Lw7cCX8DWiGV9G0D
5VWoBAcNSji/xtS7h+g6WpI0iyXOIwdDIH7fd/zDflapz2aRBUylNcFFFkwv77RmJ7xuDXiK3eGl
pmG2S7AZPWHi4tScLq43MqncxAkudu/2vMez4opuWrTmO8A0hCpG+PJHQkbF6e2Fg/u9AFcbX1Dd
XTsO3lF0hQal1k9dhY9ARdpNt9AT1HfHZAU6knhdGzQKgtTvmdSNXsKfkzwn03c3TdEWVU5uRalo
bWUXA5jv1hkNkByWesiQHuYsOD/KLWT4S5pEneeLN/ClxvlddJD+YXiyedc8M1LFL1BhDwMZ2pIw
Ti/avD+xDf/dMVObcI75X86esIa5OF21rMVajMDS0SOp+YhN+kLwIBcSZJAwqEihKiSNksF4D703
ZmbP4n8xuNhiDCYivSh/rBv0ceEys088CW5KnqNaC4UBYC9kvhX98QE9vWyX4L4tu5XMf+H/Czvu
HYchw9MghseFRb5WL0Bw5tNWx5jiX2PHdQoxztELSpvy35QczO59A73ydXZPT75RTGahDe6MVYiH
Ngd2seP3THxEzaSnNRCsiNZm3YIbB4Wv7pMOYzbaxNHlRGAbVbvqtiUYVW4OwgW6o4xeeofAlFM+
jHTqzkLNbFTx/9o/lzpuHW+kj6uaIB8CP8oQ062Gk4d1Jo+Lt3i0/zYTQQxXH6qEjGUaS7aYcW6s
I2nWJ0EdVn5ruFeGuMelu6G9h13oGiOFBHgpqaU6+qZ+ByIh0ofqNwSpxOmvxLv6fLmyYSZwDF0K
up7oPHP2sIOPry4j8qlvveQl0yQL5t5aTkrAt0Hb/VJItk6Cf6ZhXAuv5qW/IQb5Di1gUli1D05v
QRAogkd6QWkL8RAB8M8xYKYzK11plrBv2x3Z+kULSfGqyDYEWn7uajdiCi9RAnCspB29pHoTKdje
RwsP01cyu6Gg7/nM1fPvyAFES/AdFnm9EeSICMCfkNqeWAgKR/388XaOvVMD6aJQg0lhIHHieJm0
qUFOB+5a/8E6qZrf2LjdVe+LG/KRL2iPWxjIJz18zpUYIugUBd8XpBCm3PDA6hc/ZjPxTsbdzbGs
QhcdL2Nem2zsHFnk7irlpNeu2Xb0mpRI+uz5K6G0bjJ0CHfZTTBBAPpF9azLTRFBbo81CniIqnot
ezu15kjsAtdN0jIXryQ836gCUGiwaTfouSzc+vpBTELgnIx+vXw1tPR2Ya7Z/t/fDJJX74id4g1r
ogQ32RXUcl8OSaQBjcd4wa28r5UMWms0tehQtga/00eA7jRtUvN3vlcni2pzq1//ikbr0gPU7Nab
xicAz7VFEdxKq5xml/AqyWzkElwFaIuVvHrfWqpkF3pAma9JumSo9hEn7KHLnVj2PLy1wyBtEl69
7/XSjsX+c/+al9rJ+1Pv5TyYvDsBk80GB5Fb+UNB4XUrUvyFZEs5igQd38r/sjNShoCXv4MiRc/5
BBsh78aOwYxOF0YOnzKucTYhrqgAXvhGWtJtP7l+tzQRHj+2gu27SDbSj0T/B7rQTFD/hHyTlYTL
siHDrfilCQJsZ7iC+oSUUvC4i8IfyVVLFqLlUPAaUQ1WGxAK5D0nvPR1TNWiYMgjJGC2RYf15QAV
hqunq1hE/IjZuc3hkggPTb/fibL+YFX85n9/U/ZyHbnNM+GCzaJrRGh8jGBZUQvwSxDFcDWBdTWr
11gxOqLhM/gJ0TO9GbjVC7DByWyihApPzN2RMWjVnzFMieNJUsv+R+17kov48oXo5bFFgtmpYrSB
K78DPEp+wrvi56wj+paU7yU/IArc8VIqb0TKQ7kaElv6fk/coqQ/4ri3r1cJEVtKsZVFMb+rX+eg
Uwp1dmGmXa1lex+XM9YynNrPTtk3JUgCCs6RPImcyUTWvsMg5BbPDopdoy0ViiauVXaJIxwo+X80
QJu8a8M7zU2IR01nFGvsWwqPm3XF1fqgrCiFqmualljkgk9btWC+rnZKGjkAvpjf73RGxcWD915r
gcm3I3cv660NhfEvH90mzTTCxmJ1qi3yoq1qqq7O7R7IYutK6pV+jEaPRhWHad6pVnxTrAQ6rB//
nMLOpEY67xJTUWxlkWMBjzE4aYVi9lKFeJNVbIf9HP66JDq0+kEuM8qesWQf0yuRReRmTqOrMy8c
STCZStfvcItmpL+h2uyMxrS3CHoXYvrGk1s4gCSLCHWdXhEhVOoQb97nFHJNA1GpkXJzz9dH+HsV
Ddjbpj9kIvMS2teUkz9zRjW/ucoGQQTVQ9HHSgXSHxYfGiefRhXM2VOYCxYySWsiWfnyG09Lqzzs
YMNoLI/H0HwLnLlgwbGFhs98aLOMLwy96DYpcW7mgqFsdZZOy1u7jquNk+4OAWVPeHSpSqvHTQWu
wVuAhYpni6eGHllmXU9DSvwkyv/vdLWzUBUUk64zolpuEleVryUQ4Qsw8NT0Yt5rf7qPboTlGZ/n
fw5CERGkfc3qXgudP5tVT8ajnlmgFLb5MkzsJhBail5y/R/3mt2KfSmKr5uwRBs+ViUUrMiXhlmg
/Q4sI0aOo0oaq0lKj5JLf4GfHKTyuaJ9yq8yV3T00zORt3+XyGRQz4/AS0MJdC/XxyVReZkwyKbx
GIc5LQkgEJo84I8bxI27cjZC6jYq+ppHM9zGoSFqIncRFQgOxBnMQ+5bVro7UxB3OQtpFkQGFH3w
IYy39jpQ97ZkLvBPBoU1dPB8AIcvGo/+Qcrr3Ps3+K5cwFqaQn28Eby92AZCXmVA9qp9y3d7CecW
qO4SXqpjeGyyL6dFjOh2yXEgvBH3MUGAEc3Ati1J1h+h683QnzbTdBmZnA6M1hMOxAH/J2apTLVv
PIVH5sG+U1kxcO7BQv7UgnkLuggb+wsmDKEMIypOfyf3iIGwOqVlcFtYpsLB9kG0KHUUjbU8W4D8
sLWAxuoOMwaPpIRqD2eW/UGVQc6VYs1D8p8qSORb75fgp9tWtD4MIgG4vh9bg1tp5ms+zJ10d9Sq
Z6V1KYd5Agb4sDSNJQd9Rw9hR0UlSRehxrhORj8iVRVzHH3VfIvKNYNbGt7OMFqI9eerf3ib3pB5
7+YBnNLEmzq78IvsFk2nNtF+YGUr0kds7ZtWRe5esN1m75fLRIJzapuWI4l6w81FY2QUmcSAj8yy
1flXvOnLUtygWKIg42o9g7Din7CljutvceMomJu437Sy0cAKaqvk5WP5YyLjGewsGGGLulBqCR/K
HpHPfp7XA2RWnbHAW7HWAH26Py1jE+JAQiLp61j/ZPDrt3blpqyvJ1DSKnGEeUI76hw3BnBki6u7
IGepDixqxVY7JGAOKhAmg3EOF1anEYW6ElfYAjh94mccOTvCkfFJZ3OaYsjWNbvRY7M8Gv5srwUm
HRr00qZkZiwUnkztgDKI7o/zA996ElXTWKDiIWpTHj9hO1lJuOIdzna/hRCw16089z7Yd3xwsX9t
BtbF76UynQv0382SgYVobuW6jWDtjWoFp+aKnpf2kwyyYDMKanIvP5QGTTivaTCoRQ1b6A3DPxmn
0E02353uYDZCWDX3Wpw5qvV2hG6GvfJ6YvROFJGm5OxBtZlJR0RVJYQ2ZrUkXGz8T6bGKelKwnlJ
Ldxzik5+F9lDmk/TF3/zLA2wsBXm1kEoaTV+Dqicmyz59HURs0YTOmT76ROvuJWiY5/61k2Si7mQ
DGPRGP49EHENXFqhgRfXcIm6AnflftS8GwZKWvpHDfH4Jgk+MxSZYOhgNnmQT1KhSJBngHcFP1zI
yxvxCPpfEDEC5iIzS7wiugqbn+kp8wdaky4ehWoEwBG5jEDnLLBeLky0a1+Twmj5ktU5eGPaUGV0
L4QK/Uo68+KgmfiYpbFDehMtm8iBtncbpZe698sgMDyKjXRFc+M0+jS3A5mh2M5+jfmzDD+0WFLk
p+Gzk6s2wcthX6LlvEG+0OcjtLFlsn8B0Cf3XdaXxk6r7B3fGmxapcjJBiyiZx7QOFgHFyjWoy5+
Sj+/c5GS7RHFSP9eDzADR2inIYQa2FUaju8gekDMuKcBaiLUpL5j4yi0UBpxo/dz+TmFG8GT3VwX
8GY5t5SHmApqKXDM+s+BwBZ1FB7tANZXzW/SFqTaXNz351idviO5mULQkvM6omDssimTjeJdNhul
midlraCqvxLzsFrmlq5xTlPAUrpXg4WRe5pSCEwO9kOBC32wiwZtJF9lvaGKDAGcaBX97o0Yz4Oa
IobFDiPscQdjbj8k1zzhhrBBwGq9WmYfuICB4Ptd01N4qaqw6vZbquxzQpGi80dofIiR+DxlleAK
vNQm0J5iqkMY2njDwSfv1d+Zfb9ossOyqFe9rDWWFYF2lhlXCrZ7afnltr5VPPYmCzXw6I9gzv/K
VFLwb/6yTL44x5oRCYeTMdzHGfTwNr9UUoZRRIyycfC8hGckxrC+cnC5WuLyMv3ec7SQssj1cwZW
NoaBzToFheEw8Tjog9I6Di9AYWREb+Qxunl2TsCS+o+70cpRKj3GJcbnbiZxN26LzMvOgA+ElmO8
UrBrJB1ow0eok3oxX7iE8LLG7J3DjkMu/26hoHIciQVTRJxiUAGuonn6m3esyj/RB9ZJzr/C9B6w
56tXO66Ypk8ylmYLLZN8qK3yTkQrrH+eWyT5XDUy1LN1BTy0iR2LFLDeZpk9D86K8VxZbWrHkc0w
+yBfl8xTcf6glDfwj5WLUz8Zw5fEs5owNfTYcr2sd5iyIFo4+VLpzBzaM0Sy89f855VZcRluj47P
7OOLGTVIFcnyJ5vzSnraKGncN2H2j5MFwv6OXaV7cY4z9Riky2bW+i0637RAxOu2WWTS3D03DorE
MV/CGHSVMNcfYcZh8sYf/S8X2JABBk/BhV6ccec42zCpVnT7errfbLJnKgNUMyrUdomZ4/P2TYXf
KSl0pV04KSc/F4bHvrGHn8+GPhhYxS14KE5tiOooxX7t1yd5lDVkqKGLirZlQxQZ8pPYVTEKKiCm
QON69qZpc/hF+JhyDWLD0DTqn2//3meBbrBC5GuB+F6eyg8n91PTygdcsID9oAfpBDRo9VHxUGhC
AdozlRtSJmD6ajOUKUxYdROGqS6Q9bjgc2k/3XLU1yGW+HYtz0chOAHxN7RzlVZW/SN8be9PFj2/
lyXhu2w71DKJHbWyJ5EOuB7VOaD/OeFMq6GLK7fWRay61ueQ+z5/eZ9ZVByJHRDHzdfzSmVZTD1M
c8a3hzX/sUoMq510/kdBbh8CdbP+G+q0T945KEUNi25qVqIWMuLhvEYAvXVmD0OZUP8fCkATOyn/
2b1m+pg3swuAJTE0/+xM58itO0FSj7s5Niwumn1XaEsoYDu6NO2iBRA7iZKaY/2S+YqzYlBb3vD6
RBEdmo14uAQZPeS3mUSAL6wB0uxEWFroI04Ht84okwYXVwMufXWQ1hoogCFD1pPxHBAQ6ugGQB6g
jA/tqelzvHnrELsoC37qgVRC/C3z8DzCvh61Z2EXvG64q7Cm7b1s9YD9wn6XNSAGbgXImlg1agtN
aJ4R3dunVUj9v95FvIlybnwHdZ+H9pyLmrkOM/5ThNhmEwYb2tKQvcfViGpMuKfAQ+5CvkfAdXCj
tb+692UMJQnmG6PW1//nw+Bt8taz7srpE2oH/zXgIIrfWx8vcaikRUvFZEURrrGsDZPRL1fTSQrp
+0DhbEf1nL9BqR1rAgTMUZQnWlVhyveZqWZQdApTYdjSeqBOg8OfUIr2ZuZjf6hw1f5zRkQeuxzb
j8lRfmUGxV/A4NzBayzDUAqgVouaYUk//NKKLyL29OBU3LQsf8ccpk6ga2d/rRVa2vOUzttSLuEW
d24V4Tm8Idhqr8eqaDZsoPlRXez0jhcOxtupgytudaewoP2D0J1edxVwvjIcMehk6RdQd0exLWTG
zrM2yBEoIs1A/pntLEdtYG+9wNdgI0bzgU1Jbb3A+DgXV5/npziOqTrEukjASq55P1Qc6R3lpSC5
D8xISZdhu480KtSWe21erru/74rCWxET7uz8CnxSGhamZLFEP8piXjyLHPdc1UqIhPWh10iQjcUs
hooicyn8idU2oPNrRXNUwAL3z81Cowc3XTg7QrxyEiuUPz2qgNHKtg4KN4D7cUZWF6yId6haVukK
tKb/369jEqHs0yV2/45cZb+OeCEDo/xclGraRN7cRR9frytklWyW+T3p+uXDCZp1PP3+aTzjaHxz
PihvcM9pi2SiFiyj8jf6jYY9HFkEm/sxwDBLjBWhCNrSVu4EF9h/V0FIiTs9VE3mvxvf+gHTzl/a
rbI0fkVL/bNaFTLiA1c/T0mTYJoiQrFRx2eKU38QY99YsBNzo4NGKW6ZmFjGgBC1kBz0SXADYyyh
dktneazn2kABuQniL8HWIM7GK5itBjn9SdZZAHKCRoXrPqN1VEtQoBCBz4YCijv5c5EGd8ukAEOx
P4qHwPQRzcvPCUxSR9pRDgNjZaTSUnYQ3uh6lFVG6IYbfbY6LzTXl1xH2LfpKZbm9gVuMoyIt6Ay
QJr7FKUTklyLwMCd+qv7mALHpSkRyd6c2kt8IQMnsUt5/G5niKOmGtKwAG6KqQJukyQTbcOua+zt
G0UoogRyLPYKV1bxpObAob/EuAS28LFeELclBwk8KCQ4CafVOzDbC+VWn5dpwtxDyG2MzouoLN8h
wi+/VSZKApJOL6bYymBt+zfpI9iVeSI5y5q8t4o03PoHuPF7K7kYQ26w2IKRFiBGVfMzVBGfj+/4
+FOp5RC354VsiOzH/z0As1dv0EBuwgwBF/B99EIIZDeTQCOcx1Cu+cTAdtIJYgXYeL+CdTDlPA4g
QurOXDLgpF5pNo308v1xtmAnqcudauOOMTZ9EFMiJLYxE7Kgho6QhmR//YpAiJL5N3zfrJfFUfwQ
xq+GLZ0oGk1k4Rr9EyV7bibKmA3aoTBjhkV8/BBjKAq+/BVJQeby0Pi/SOiHysl9OhvM1EWaJHpl
IJSCVN1carQ7J70iuvse2b9gwHweEY2E9OhRCpUrVuo+LRhwckiqT9h0zviPfhh6olEK89Hw1oB5
KwM7uZH2RKRkImaZJOmKr/uPbQrmCpFO58oxlP1IfvJOkk4Dy4aF8LKFPhzYI+T4O4k3fvVBFhqE
nyMvuMM+zoDjliJ0PXMRMyuIri4/YZhn+czFZPVUik1t/SNRdZxaP2kkqB3w7O0sKxun99HMuGnY
o818+UwjCo1x3bmlpjoR3Y/EXyjuwMLRL1kNzcoj7/jV2HflE6GTPrwGzQLtmFF64deO8cJpHbVq
coP8/XsSeJPwGh9D46nsKTUS/qESasvbqtWLFKSNiWHUhhisDECtb6SVcYtBxYXchrh65uFf0Mgw
tJDU+v40V8AGnWnLmkkZG3nv4OSsm+X43FFgnvy+OkUUMCzLeBfMq1RDe1WHIz6yKTigqbjzGMRh
oHdMRfitROltp4u5+puQWRHER84haBjNGuA0xHzz4rjGpE/iwh0UeBXA9eSXPoxW6JJnNjJHzhXw
JAobsXRrzRl2tG7qz9WVQD+HzkJwshMql5nYt+zL4yzDuMXH6sSQg2hqO69T448X7LBHtLqlhv+/
RFPwZzQ908QFOYvMCR3YF8vwx2nxWmh5JIsy0lObkwyT3J+lqO8DMiJmpPm7UHgTGYVVi7tivTYG
wafxR4izzFBpdB392CPJ7gVxOduqUHCz4QoQLviw8Hxl44oDLbuHm/ti5dW0zeJGai+sjeFTVCgA
PmECivgp4s/OEZI0UfOCHOXLMcphgGWxu9I7cRkTO+WnhFllhCIVhDcLcmxOxe2qTYBW+8QBMNVu
svo/U9r5iAUOx30wAFjPUxYiR9ys0Z+Mqe8/Pvn1wrpirnXrdU8REpSQS/PaGKo1A5zHsDB1e2bY
/Cq2Vo0Nl1dD2WTantwi/HFtDCtMpxT9PumZGYWbuv4C580MU9ohYLq3fYKd6pY3rlIzUG2by/lj
HEA9p9whKqfg+lYXWXscEpwCkzrvPDrhtSHkeBONeSZc56un6c3Bs0PmSj1OgSrKpG08I2y9yx7a
geQsaq6lMAXqn+y5uPlD0/6teRihJ5FPrDtvauV4nKPQ87IMS6OOHeOndbu6r6jpghYTP4et8xRW
vIvmcu8tPfu574I210y9ucLjIfowmV/AcYIHVrsd53S99m6dstfPG2WDTODflPBuQQDAE0obPzQN
7q5q4r05jnqRctQ8nyeyQkBDiEdjNiwdtE+r5rR2g+9XJRaGqyE8HYqxJh+rTeMh4uZDKmD96+po
JxmACI7Devz14CFALrnHysSsgpsNgMpZSuUUX00rNFrOipoovE+0MC0Bp2fYKnPLABp2vXjIudX+
otgg0jZf23NJtgKT1aOH6F7ZVnkTm9njWCBTDcG2gVZ2VroHi9t3WiTntGnDGdHjXhO/DaGcrLwi
le8kRyjZVx2nMwD22mFPjbvFey9VWPo0+MlP27sPzfbw3ECgDrTLXEscrrnyltG8L0AlFgMbGM3B
J1QVyW3A/U4Yjk0S9Jg8sK3uEoQk1d4hVs2kXQOt61hNZ22rza3gvL8VOTPLznqDokbDvxdeYwr/
SUar4wqc1MQD6FvXJqD9xcxT3I9UW/hLShPTgY/lyh5jYcVg+CMQo5TLJfpT66LiocppqUfASm87
wlSP9xZaDcErz8wOIcE+LvNk4WkFSOPd31OE4+dCSE57Y9XxnPskQ6qbKoNItFywTCoWyJHTMOoF
lVVYXnQ/Fg4DGXXQyedC9i3KxllUKeZsTURjdV7uyyhDY2v9PcZYnMKZSPQNsLJXqglHgFQZkb74
ENDyeXL7LufSwv64ABa0R+LEh8EtlReyR8rhWE4FjMb18YZv1WsTnbrCnpy9fdOUZc1nNM0XAxc7
hl0OliTYysOD6U/7H1/ZfQIovJvRw67QsUcfEPw62yMyJMQVJHtizfmM7bd682BzmnpRpR+zvnOm
0gzBV3VHQ7ef+a7AdsAefPYLQxGEOZEiTRhlGF98ZrmeZ50Qt/IKxiA56YopWExNVmgSKYu3qCxI
kKqnCjAir3EZkiEMpqBJIbVpjyv7hhqc3dRRjoxHbjZjoeYum/4HMRKKyg3U0GmQf6RC7EVOa4ie
va2hbX6O+WL7Od7NvmCcazthMfsqNt1+ZhKl6mr4yHvwnDzSwRN6oKJrpdGYRhxyQCBya7JUe5ZZ
KySVgYiOqdB4V/cvPMBdCIBabJySfgc731QQUHjKPf24CASCxCFnxQfs6p/YWbYOTpLSWrxJ+G2t
J9kIyxNC8DgVMrfM6uNfnyUNdX4IrwPnNIKhbk+tbHNqFz1VMq6SXKp+847yOqEpLCDyhEBSG/Ot
yni71L7OI/LLfYB3pbadknxeS4XwFVQfr20Jmdg4xaT7flxGEApJKNHdpFvwcPG1BjM/A0zDX/P3
b8wZoSrteTc5ZwkelaWyCN5hNxUI1vqgNVAast2dMlFfh0lmByOOkyA7EXXegtEPvwONTAirmzjh
xY/lE1iY2WlWLzszgmDZ6nkEZcY7mkIYsIfMHnG6/i9MEpyjIxCn/KZeV5kHd2h4PFh87pJm314W
DTsnv16/8a/TDonO1ijCTl9FluGxTlIW+8F/p6LLSJm+2Pv+OYaP37WaWBYwJMKJU4DGKM2HVyIK
AQHZgr48P/NEB4cSKL5XskavVYBuuffdaU8q6OLuPbJQiRMl2ydsQ65oHMFK8CZUbLAt02rcQrtv
gLtboGgtIW1VMxpMmE5nnAA/X65bt/SbUv4AZEf7xmdmPq5RhEvmSf7EiBgnzYBiUZOwixkWSr17
RfJpH520LNB9Yx8OTfKN/LbWkdxeq4LUoRInueR3ZEkeeSC6TplfxSyg0wTpQuO5kaw5SI6RXWmZ
nwRLxjuWROkeEqwsMnDRtFHfvmYY+D5MdmSyPmrYMSuDefwOIhxAdZMB4vwUra9x9OEkl7Dlnu05
xKHlj/0Eahrj/RNfXN5g5R+kJ/ERizt2qrhByueNY/G1ZDMhhs4oi5ymm6N0COziRVdPrYqfTbL0
IvB6kXeXJZ9Ge6OteyKEEyDmHs3KyDTzDFiCknVz9HHtby3gr8btxK/RqwdM5I4EpLFYD/Xlbr5M
ZF+245jGHw/WPyiLpZFKzrkvwyDWYN+Plpm0gmVlvLLCZrTv1ntSReW45S8AkkvjHokUyLnX0inO
PcYbYKJMifos/4XfTj9A3qyRFkDt/EXYkFnVtezLjsJS9vOpFAHiqd9FfQz93PcUl5gcnLwF49UJ
58mqrZPs+kWASyxtuR3vPs7NiUtHvvhO9d+kTDKowfSatZkN3Rv6rMbMWCLEHHgs6fXtW/g9mY6L
w6nOiRmuf9XdWrexHAaz5ItI6Tdc5Daz4LG49hP92NjhI+LlMe1u0c/9mOvcwr89acPgmxh1sD3y
3nlGf2tfvwfUb/FPegqcyxMLPfGLCdgnjJYAlQnfMcl/XzVaxUoEqglTNTFjS6ymaUXPF8KKiMow
ew9uozc3MskVHQWvU5qQcKazQ5cK0wMPkT4bCnjqdRBjZQcZMAAcREaEqcNERpMSjfhLcV8wKONk
naTObd8VVT+mk0TSYrmWHOUErNq0kt+EG1Y8rMsQwXE4zsHTvb2L8KokjWv/4akEZq5Bwk1fZs1T
kyN5H87cQ2AgygRvw411Ts5Z9C/ve2NT2gwH86e6WDtu2Fz0HjjigsFeaHIkC1NyyOCXSsqX2RkN
7ETA41ue0zOS4KHMVVpVUzOPmkjGk7qpPeOajarDX8pP+4h3o41MS8i2HGnBIqxbmIXEgCxh8IEs
PrjvN1g+221jTSqKj7+XOdC3B8t7AY4drbF2vbjAeEnUOqkzzi1uix8wCE/cJTdoxFA3HmLe6c/c
gIVSEpvjEUSHhYAs8PxDyTd9nt6eJHrCo3aJ48kbMJfTT7nv7e0edHyP1uwRz24FuNO1QTK7FAF2
0hA13nhLBUjuwEZDDNjfMUknlOAQ3FZ0u+dK/HwYsEtlhSMsOEGXfkVLWSwNFb+nGA5JeWq03sEa
gSHpjize0I7+vD4pnLhBrkZdLXSJeKiafHGe7B/mOOQ/YvSuytrKnCFmSumWyPaoahuBVubcM33f
E+ETp8y0bIinjcFsNV3G/0DIAZyJJDhsXvCNkW0QZAoGJ/idRJNfklr0rl8gEtbLXkY/+OQigp0d
mbgEJySgCoOynv30hqtsmIKB5/cup/n/fhXAuWH2pqP1UWz7riS8b73wEDGAn+1MfMJg6C8EPH2C
braJrvTYTqgV0sG3LN0ZtpJwR51/b96ZeMl87w7D+zl1D5FTdSN7i8YWONK/ybwD4uHKWeGxsDmI
eBk0P06nWXsv2tBEDOtrNjio68L9lPRgqsaoyAhJtRbqYtO6jw+nNndDPKXQ8r4Eo4hAeghq89ot
3fVFknk+rCxVhST7H77IUrIsPdXTr8fCHWNh9WgljH/WLMAX5NiG7ZJNhwUp0UvwihvKBjLzzF+E
6e1z0agFuj3BYsZKi/qp+5rAtxCGvo/JOdcHhwbvFi0U79OQXLzLaGKQENtw6FoPXYi6VfyViEOs
GXhhNljpB8rckYwEYE6tCLjKlPLzSv2LR8NnUXDfeSY3hPjYEGa/1EKTXoyVn3pXUeAmw/6f/DmW
x4/c3qSWvPOxgBNEZ0WtvIH8u+1av8Wz9AIUPsneMh0Q1vh5AiwLALqJMTTC3lUnOK3Zw80SDK4F
LBcurpQNFMSR6kFCu06Ywdat86Eo7zR9Hg66Dp/6ObGSBJbA90MnmqmYIy22NwpQdginnXaD4nq+
oEL7JwTo3v7nBP3QIKFQHz2yFKAdJzWDjJz/cwidknyex6c6dx6WOjnqNGsADei2CK82cNYYrG3J
EnxBCOqbzmgp0AXmwg8GUe3lf5pb4Yl2pu/9D5m/uNLJ2DLDSHl8d96VhGzf7iUnPDqtYOHqeA8q
0E9/enuXY3q/KeruRzHyk4bC8qr0JONn4MjdaB8V3r3VTmOT4XAVgKs7jG88n84XYWdILlniE+0K
SEimHNZ8zBO72Kj3oeSbMjv3WxtoR/KvL4hOe8WVIa8b1Agfzv9i5Cam4bYatEoVFDLQl+jFXSL9
yWWCPACH+CTIihejF9AmnRgi1clFOIiIY8XPQsM4fVT3n0IN+UUpr6owAfvdHqcNGeFlzEK+hmA4
tbklVXlllb5M+EaVRz86Qm7kzjDoMCWN8dHbK5+qcI8Yjy4L8CUa/rcXcQXurwnulbPgrWZyCr8x
jEzwAIeFB1cfRPAIAbFuG9+1VK4qlBiiF/TWiG9yvkjzqoYe8udsRwYKK5hSYwYG3Zbp09JrjNJb
3HAkGuAXTHt4v9pec9Y8dCK2yya+4855gZSBD+7mkTyRqx6xppKQ1L1xuwvN5HSOdpGXqxmzHsgG
8Nmm5twlLNcYURwwDZjXA079SHbgRn/05nf2T77e021WdVVFVbh8GUecE6g+26feSkJ+5gqg9B1e
JQNvDH46LUbRH5Yvs0ymdmwvB4kz8Myx7XmFgmC5flnXFGWIqDQEA+o9udl9IKkQA9Dye1HBVR47
/NcbaE5gkU5cFmhrJT9uIW92o67U2YXn1HSwx3gNGuDPWR3CVXyrdv2Og//TD7hyaKdrQCnzI1sM
8+LPdQYWXtyIohgcW7v8cpk407UVlN3YzO+OlTfTzFOkIYoBcwQ1Z5bcWsSYPSy5noZmOEU8A7ym
MfPPleJIUEzvjTkMHqhBZrutiKWoU1XciCS/TLI+UMVA1dhZuT3TSVDfg/N9fjUIQsdpbZMkIr/n
TXLdlq5otTOq/G/k4QIf7M2k1k5mBo+KHmoIBNj2CL1tuK3bymw27yf9aimdwI9PyThQ5kvEVtbX
YRKgGO2s2Vgssbx8G93dRlAkk1waTi7mb+dLkG7iKizhzUjUZQ/JUUI6JNnxcGzZmi8obXR/CCwS
Xg8KpCPMxcakawf6Szy7XQcdleJl3yrOrv65hBYNdRbQ8323POhn2JUlwCZ4ElkRsHXV/JMX/+6n
A0Wu4WLMEP/A69+5vtn809C/OvoRtiGQOK0N0t8s3f3l0khBXMSPeTYFVVrOVc383+rqkTq3jLOL
PQviuaf5EoY6hWNjAQ5odEn2zP6i+Ij6nXNja0bFEhZ0/4uQm1PW/eIBImQexzNdfHv79VCQWIi3
kb94PFM08JGMhxd0+PsNoKVRTzyJROoeHdCE/COvgPiK5C7U4yBYhwTjVW6DhWWsbKkOTAxiLiAY
8RbzN/V5bK0Tp8BgA4wnqxUSFfxz5bpMg3TiKwRvT2l4WK1HbLrYAwRe6ZCiFWVJxxIIJHHvLdtz
9iLrfsNYczh80CrPWlrazdjkAlUy5CgsE+rLXpyWf+CWC7AIHV70R3pK5BaeHWgVlkev8B3xV85J
B3M7J0CSUosBj70GxqAN+Sl4/DWc/LWDIbvlzZIpzZ8b3Ec3lthJ7C7/GKJh/ZwchO0YAKlBQwgK
CO9ZtvUj9KZRO36os848tyT/nRbz/zEvMRqUOvi/Z6JLo0l7GnnvgQIDJ8Q0pHIXs75Ln38Cx+kn
3YpmJwnyyrps/3H4Lm4jTUoPfF3pMOnUQnw+E1zeO5vSa8F7M6FU30pKz0Zsg5ui0GqvFnJqyyS8
fERoJn0/N+jDNz0xyb/57CxW52N/mjcU3uKgqhe66SeDa0rH8Qdk69hKpTd9woVj7074K3iD5kPp
wRskKzzEz+7c12ErUCC2J4RhgPg9yu1k2X5v3LIzIgkb9LiuA1vmuEY7NzYsY/0Ea0RDH0roJTkj
wPGLgrU5i/VZWA+GaPPap4lTNWUoej+Zg4fMzhkFo5mMeyJ8cSMbUUe0Oi9liTaa69lgA9oUzs/I
vJtxCc10uLWUs+ILtVZT6aa8+Pdj3J6qzUu8vvMNMEnWe4T4bs7OcYiahe9fR5A8lY4yqbmPU3hp
bUNNercXHUQgh0Z1vryjiKf9LQMC2p2q8kvyKu2Nj4MQK6yztHca+bRVKXHEscZjcNYE8R3GwQGh
NHkRpDW676PjKut4gmjxi4nC9qf6FToiV4/0sjOrJX9+vA/QYlmaiUPZRj37M1pA49IK+ILKbC6n
+TBaOObsDuhZkOgLofCqPfmE7gw1h9mG+lWDMXWCBiZ0ddIWwKhixNv+7qfiabDxoYn7CxOBems1
31BHlw+B76q3CkBfim7iqNFzt1+XZtNEtq0vRhLnftjScFZnKn8bnJI2pk//bkwVGr4lcmz7+UrP
D2xjtN/Wke898f6tYE59ynnCw+n6zm9ItWLh6aXkQOmCe0St5yePTZlRVRW6+/xDoQJ/B1/IVvhD
5HS/oWrhRgX8R03LqYMqI5mOJUWEuoiPL7N2dMNmNOHrmghvhMXcVmZ79bj/u1tn2OP+b7Bw4mRL
DgKtJzx566PPZDZIzD4T5AKT3CkiNBqup7LzI4Pms3pk5MPzLGGCATap8comBxLz3OHNMAIQVCQo
tznMxsDTZO/IGeD4fWICrlTnfzF/Om5RxhmU7ct63QaxuVOHqih3krJ4DmE+9cRy4LrF9YEpqK0i
bQHheY5AgWOYUEGJmaK/ZrYYxC6OVlu7znJjMuuL+umDi0eKQXpxwyn4/5q8v0IsC4YXtt3Q7QV3
BhRf2yeTmQSWQKZftdyxHtNjscVpaatJVUCw5tX3CoNFLC9zJWuYbYgferH4xikwfF1IsGIXxvYo
/kAPU8DH4mCBs0RWig721S5Nn0kuMTqm0pnVAYXqr5awuwZPcL06pxhtdsntT4oxZVnb917JY4cf
WIuKuZ2Sz75JplKOru2tAAesWqe+rlGjLMXJj51eDpQR8kaFW3OVWrFsd3NZob7NdbsFpL9/S8iV
idEblKZNbgeqmJ5FBjQFX3h3EtVHPy76XPGPIscMChwRMg4Fff8k/cT9821EpUI4uaMWP4JHn6yc
N3maMu1iak/W7JtnF7g4Itf1+UoXpgzVnGhiPck2QpS+cZid0BD/i1KtEOS2Q13FL26Su+EHpXsX
SV/xsOZ5eN4o8NsjBZZdlEKfpXmWX5qjeXFOl3I+lOSMHcVjUSPRXii9RQ16ZX440kaFiDzQgtvA
PjOYBMJY+5/ZPdMp9WA9yj9EuoGTR2+Bcz0tMJo4BDJuPAkdh32OA88+n7lyhkrDKNESHEEF/DA5
v50nxLBj4tIr+p87bAOqr251zLClfpTHZJs2PYAZWHIqcUYT1ddwxYjo2kgYIPOVEccYKhmIDBtG
rZrz3j4X+cT9cpTjHne11qlPsWCodUMd9tm/6maLWpg6l4ToGw5Ye04zq+7NQSInAmvSwNtOrlt6
ld4mXljWFGU6gC/zw8+HlZ3FOm/0WpKHzkVDTomCr9XudrIZ6/LzUTGQmeccTpYq0wp/S9/oOuO/
nOOfxOTdGPyO/6fAsyh44NX5hhzlyQWCRCjRvF9Wg/pBlc0C/L/aTUDvX65FuQQHxSWctWarpULt
NqRju+AM10U/jLNX//JGgkw4pIMRJD//tU8zfnc4e9RsuMhJkeqQaAmaRsnWUwsNA13N1v4lL+ha
Ps8BLY+B2+DJFTOSAp15aPyYbRXBrObk9m5ZWvgcJFLTERgKn27I0OSRR6Qxdd3LpcEltRWmNyP4
5os7xRJ1f0ANArA6HSDDdLwM3xoDKsCZLY7ChDqYfRrpPdn5T8MC0cWm1fBgZSK8CrGuufYfz/Im
9LzbQ6proPG2zSQEEq9TdPUKrGUH+/e7voKsACKNfRGGjf03HXx7zljCbQ6GDUyIyBZLjbe02mrq
nmIA6jN1nfi7Xdy9KsbgV/ZUt7GhLfsVdOJHkow6uWdPEK4cfPy9LhHD1EaOxk24lnlZFhCr3k3m
U/0tsFh1pdDk5CrRYJ5V4YEOk9EW1i4lC0eEJFcN6NhOCjoSknsJdC1iA7/aVGEooQZR532WxZkM
c9ZFsWuNEKqC1NC5Frawio6anv+T0P0Mx8gXHzovB/qwIBoWHoWzyMe41Qxlk0cdzVtC3OEV8HGE
XTRg3ukWWUi/WZH7lL7yyw9J47m+Y0f7v7LtjyX7d4hfDVGO1CwBGH0Xz4KcmMzeKZDe6YDup+Fj
PK8Tic4g2yatMajxyjy8ftVmzcH+rUBySmN1UUWUprgkNxaJPptgBepIXLYkv134CEyk0yt/iWee
nQUukjQ7RXnRxYqKL1NjoaoTQEoVcdzqFENRHuijkCcy9UjEM7h8BFFnT+6gco6ZI4j+7DYVrl83
ELQOSHGv2DMDY51PFN5MPzmHWTbmWdJLZuqTJnqJtOofb0cVDsQmzviD71G+iC6Y72MNmbKyQv56
Ojf57sB5cq4qZqXX0/v2/ubMsqiGAWBsCSD6+He7ev6F00s0ILeUpaPqmKkpkHdAYK3uh5vn51vb
c2GPnc5nutPBBX2gMTL20EyD2EceqVltCgFLWrmNAjM4zbpArT0TAkkPZs5eWh00Izahwfe4Fs8u
pKOGZOrRR1ds1e8XZ7sSjOB1qeKSNGANVySjMT4j9V2r7+XQD9j/znxf6JKig09Cztc+XJzTYHoE
m2wIgeKEorG+4f17zJrBKj2HGyw5Ja3RscIjN4gs1iDt0m8HEieDrRDNweO5L7TPt8OU/s5d9E97
zIX8xIBvgkS0qIFXn79BeG4M2g3ryZK+dgAfu/khCwyqYOopLu1/E5iJWRkt2THHK8/2AhmaCjss
+4uPSTyGGSNa++lPzm6GxO6guj7wx+HW0lkH+l7SJHKkjetC2BAp59phKFCxI4Yr5rf/KfOLRQ7M
2FYILue2n3TLda5qB/U7Vc5TlWk+DH2jKRA9uJFbY2eUZ/iAyuc5AXVHRw7913uxIhGG0f161ES6
UmRF9dkqrr5WSdZ8OmSX+nRGz4IEoKGot8P1oyGNzcqTNrLB09tkO19wy4Kc64NYL4VNmMzZLixr
nYE5gC2/geMbIaG84PidmrGYQrP9kYKVPI7AhS4Q2Rnu2PRQBYICvTJZcSBz79BLOuWJ+H/VR2gr
Gvn4f98P7qccNN7nXVKe01Fa/Z3ZarlfJoP5aP3qi/UEajbvgC98G+Aqr+xkMUBc3TUbTb7Ky0x8
0cg7lKu33ZLZpcYe5cEQaaZfaAedVCeG+MaKpoxNRXneBRAlPZQp18B99HAFlNW05cVMiNnFgaO1
aDBLwEwBRFi1ZQEOolhmShNCQnaU+xEwScJRmEJnSUbbgfPOPV/sm/HSR2on3qBt1DWZ5E5mQOPv
C3RSoaKKjxds8XRnALAH9XzGMrPyvajyGOTbhMTRpAafQwdNmxaZ3WFYPz+CCLFM9b28ywNnOMpX
KpBASVlJC/2LoeZAXkUBRk030dL95iv9nk6EEgz+r8lMDBOIepQw37KiIW2w5UXzDUrKSbyP/cYY
Fbk+4rfuLE6LvJWuFKyRGI7w7V7HWLMi04VW988RltuRpN0waTm8fJsBHuYlB08gQyAUlhlHWMJF
+iMRLXibP0SLGWIVhm4QiTcYbsxiAXdGIe35xmqTj+9pv078Il8lnvST/uOjWGauyuuP4CBTfPcx
hTk1Es5VOayMoI/xmCa2LliCymM/eLPNy38tlofZFfA/J1vio9JJHQ7FEQQJ1/BQcTU+z+KW3qwj
vkr9RwKcVMEl2r9dlTj/bow+916g28Vik3yor4pl7uHlIx2sv02iK+cRqGgUM76p2oDhzpzkonTQ
IbaV9UWi88GRHcke+S6h6yrszU6jXQLui39CRij2JgTF8/4OixWJrJePo6Q6uSLP0Gu07byu2vq7
IEZgIDPd1fu/TrrGfUQzMpnB6wBYjtgLURwdHhtKOBXIBaOv1D4zICTEB+yoz+hRNPBlNK7wLtAB
CQTVXW8Buj5X+cvU16NMafZlVN5zVsnYOpxitRCpjnlUHuS20sS1zkO70XJ5DQsS4Yfom0VHZbe+
lI6gnluFUCLKzCtkd7opQoieCqvwZ82dFI0Rtc+oh6lxEYnr20MlkSSoxGbYFW8V706laCYUf9dV
b4o42SiR72K+NlLh+eTodQdFdcKs1o9IoYX2FpFFoxczHkjk9veXTR4JgyEibLN4BvU+jqNQ2/zi
H4cqfr7O7leFnF8RL7aj4Acl8C0tFbKmHZKH0pFha3t36CjkxlthI/whHiMDsm+RsgaNPJLJ31Y1
y2J9NDhZ5FACDdiMryZZwdfdl+ThAOk5RjKxSuiHvoQfn2K1pC7/VlJBNE2W6KuhI6gbRB8VTgZR
rmu0vQ+LU9xCAUOfRX5MgvCDDaMD5bPXBViN2gwsgaS0r2QGQPqSeqKWxnSjQ6K1ApV1ntTVR7hV
gJgUqxF4+jzGh5SXnZhy32BFoBGQwnBG6bbrQFsTb5CyXF2OVYCHRznRMu0jFgiYBdYjKlplOB9h
bhfB/Yt+vhb3fo/o//IH7f3y9qnyp2odJgaWwI2K9qUhdBc0lArBTMBmIKE6J1DOyci5AWUnoaUI
FgTAtBpYeYLzvrXBHxwP954ewY1ErwzKmCG3vxSG7RAQnbHWeH9PrRbzwgX15Sb0wRjLXXXJbCbn
0JDqnoMmdUQZqHhgl18UN1gvLpmNXsxLFQr6EKcPGpmaiNUgx58AhWeKLMdTKbYbSZ5O0nJxwd9K
MAdCvodyAhJg6yFhMv6IU0x/ce+j+TSzsz57pNKND6tPww//+IB2mZKHg25Q56EbCH9poeXu4eqm
QHfQCqTx6CI1ItzZlwIFyhlnHRhcHa4mCNavHE1DhNkc+CFKr0BCcZBPy7tIBTiYipewLX4oxNEe
kGNZSo9ShuTf3sJzHgxcsCWinarcmKfsTHVTg1SbBrk2m2MoDtR61OBndKjhnugHuj0AbJPFJbCi
vXA2RoDhqPvx14pizAmW0n0MA5G4v3VYjYJBbo8oCTWgQ++y3lD9+KlTNngfCWE3bubQkd5lwU5X
HjNzp8C+dIl6iuLpQGzgGIJX571ir7+01s8RNxLjVhC87yUGOFcGXi/i2vUSftmcrY0oDDOGgYXg
0jZbSJo71jGrbDeNIr81p2f//KW9iykCR86UBgdamEvcfgN83JlYM/7ygBIgCYktajig7wTq6zwv
FLwwQjKNFExG9S3ygJc2P/gYHMN4+a8x1G3ntSq4sjE/BJopr3LMR1g8zHi40ciq/ZLG7a6gV5sZ
6veaS+u8mHmHexxsR/hGwXsS+3Mq0HXvURkzBPfM7wtHzNNLaJXV0T61hXKJ6JSkPzg8IrOR/9fX
O10U74PjrTuAVI6uoNF3m2n5YZrF10cpqk7/whK4Mx1qQxwTy//E6w+ZZ7MeX9GQtUksILE1N7ek
1dTfVOj7XKwrwAqadk9jHWa7Q24t8oINM75ixS+nNvW+9TZWTVeMadh7TEjgy/L3tM+2RHjAyn9b
iqpHvzf44S6puTrtho/kWDoMFEwwNnBReUB4BSUhd2SmRcrYIO4TBy4ugE4oMEG5WoFdyAFZsEqR
fYwrfomNJt5ufIYOlWw22RJTs45u+IOIdvQ/Cjm5he2rsq2SDh4hB4bnrrVymaExSCDXUBHPKxgf
wyRf3oxA6Uq7DhQpxeqeFVjIrpEishak82ceex8B3Tr71DWsLWwMt5L7gaEP7FrSYmAdl83pS7lD
S8FBob39kGhs6LN2gdcEvpbuuwgV7PTzCyx5eDZlJi9UDk7jsmmHDJwOJZkKu837IbxKLtcg4uoP
9TyWDCvxt9DSKJi6iR+gqVD+cz7+09LOr/RFPPF+coOmOhLYmvZ62oRFkGsFBCXsk0hJdn8XANGz
cfRAqTS7qlW1tsAFWUDYXfJbYfhcWr+XDkcAwsH76yxmUlSoFsKQssuYrWbiEl8NDAQbhKmkmnAq
T1y2RATc4aAd0T5qE5q0Teh0bsAXl6pz+RtcGNp0l0rqKpVxyNgipalCH4VsPyF3eCa5FNUxTC8V
vZGL8AbTSne55lnhUecJvq+8amlwZ1gyD7xyZt+t4cizh/1Klo2gZBdak/LVV5JfyPF25SgOwAqh
QkcKvG/flOnJvB9s0JKtRhr/pqw0yuM9UXdayvYc3lTZTpa1pyWqoaUxP+jD1ZpUnUKiOsHrQjrp
Q2mmlhURLKYYnOly6jX0FnGEM0ciEE4WEkuF2LWkm9WjgEfdPCIGoiDjH/4mPYD48GXI1FXpv3If
ShcoTE+WSW92U6+vvrUu8C0yzkB0WxWQoHGv5urpzDY9gR0/83KJdL9F1sFAXc+3KODiMdpikAjo
jQVuqkVtpYXL4GJfQJ6ndzPBZcUQIrl+ce6OWJ/rwj1XiVgihOtXGI90QcszPsBjGIjK0m8ML6Qu
OLPpiaZ7kLQmlAFPGVVzZQHIXhilsijL0mHD4/N/3qQ8ovtHT+MTtT4byZC93J4qp3LJs8HaZTOM
fyoipsVAJu5KE3d0jWXl5cU/PXCfnoUAy/dxvtpJ7BnjbL6tRQk8HSLWSE7W34WcwMd2H0eI3JNY
U5erTjpYeWzg1XUWeMvVHYppaLf4Om+b71Wdv9mDwM4924z22th69wAber5RwhGGFjVryJFRlqFX
4jVzQWEqAGZHfQv3oxv9C5eKcTPE9xBxSl3PsR/Bcx3I9Ifuikd1nfp42ZZ/tuezHL4N8J6lVevd
N0COJtulKQr7HNEoxUE7doJf35no3kVWZLS1xHXXhIkCME90wWzbg5XDl5nIEfi8TrwlmXEIgmGH
QzfUh0BdU1FKbwRTVcmsrma8FMVmNqcNah19tcAZxEyrIKPRQQbYHcrCFjTy5jD7lmuZZObKVRDa
5Tv5c/gORg/ldzO36XF7yp7Uzfi5tOIjGkBHKou31SAp4Jmf5arvuqlzX9jVhCViaDiyPyUK++1X
RAKAozKJwm7aqSEnaNF+qbi8Y67n78CRzNCaHaVILSDLga16TQLC8XhBsuhZkNcm/xftrTKYZ8+Z
YKgJGqhmRS1ljn8dRU9B5WVEDuKHvLRoOm5VLGhHpe80ZhesAVYGBWjO0v4HS5irGGkgGXLVyfLe
ny13rcqRV/F5QcDjWQJNMWpK4i1zhlNWSIIthpMGhQadqTOQ0+8/01RBO+PLIjet7iaAIDeabzFn
FWnPTqi9mlqVdx51JpnBAHLmxqjBdTIZENKTeHHMqfWPeQ2HUV1u0M5V56KEXXTViUbevgkle0n0
+ypmnnUjmlNs2gMexrv37Zrb9zFLAjSWVDdA85J8mF7fU3sqlz9FrTzoibV66y1OjF150M8eeoCB
TnUmtV95K06uNlemUNTvPmIx212ojOqwa7tHjnydf1UXSlvlTgjpCtj/DL6WffoshfzJ9bnlq9Gv
SRaVJ0NsTtepx/u6gqdeOKPleHwL3xeJpqebyuSmEMkqLy53MHbBr5zqFdtcZUHHWjlJ+Ya/h0fq
b4HJ0kpeTppqqTYOvSI5qyZ8zUBn/tNLBrhXjXsSSNpb/VDR73GWod5+Pa1MUXOwlyioaFHDYEyo
enXr9GOk+RK/EBR1cX2pVwheVW/LlaB3Ov0TegZ8EHYjKB36KRJjUT/MIuvyxTo9K87f7JatUWtT
z13JPAGKfuaU5U0jU70+YVEQWNRaZXRkcFhZS1ripg0jl3N3D0dqusvHyEjrapb93qSiBHOQWyxQ
436cInY5t4DO1q+mchdjuNY9ZRuEjiF47hDLNMWGv/NIFTMhTSIq4QDQAgNucihPL+nLSJx2e45w
6im/uBjR1D6jeAyxaedggqX9f8dZsFXneIVWiGULzBspgLZa6NELRBAffoK2ZBcrm9Ut/IPaLX+L
XEydWLB+KfgmPJ37yAfoGpcA/P8Dw2LeNOKGtaQnQOPWBjPg3vlWJeezixqlYqtkVh07aNbaLzaL
tQTzPL6udAdDR5zzMqVpNCk+D+E+nx99PfRAgWnZ2Vs3wZVwG+g38JZ20rZw8CisjswHU7TS9Bvr
iLi/YoTQnT+4j3SXBNZYeIGjIKc43nMohgeY78DohbNjiJ4OgDLEHuOG3/NdVE3RJqmSgyjRYrRE
uMuOht0ni9LfM83piq/NGuC/wxtM47fTyVdgpkjlZ+zOHYad9yQdQ5cdQ3izSS9CC5xsk1HlsnDx
mcf4JHdWD5sGawSq/X24HrFMU/CoJ5JVuevJ9Rr6Db1CTV2BPwNxHqtFfAWYjc3Ajgk9ncjW3uNP
ggrKgH8aZ6GaapNb3SJkskq5HdWCPvOcUNmegWYxQHAZbb652uwecZ+1wHzvjyM6FOCXrURB6Fn3
KCuhtnYyASzdf9EQ99e4F3F4IsBpEn+CmGh8Dr3g5TeKB/rGVPuqDF2lS/A+8N4TgsHfwuXdIkvb
feHAKDNyH6+yyZKC4LpETZIZzo4WJT5S/AlYDrEZo5qbxsXqXUPe65Lu6hMp8uiYMgq4iO4H+IH5
SULNWdyj0LdrDn/4J1fJbA2HFdclk80H8+puKW+ymWCFkgOCONlL0M8h3q+CVuS43rMSZozO6aWE
9vIur8NFmOOON0+hKKSnS2x9tOVDzKFFmbaHAqnWJyfQh9f/uW+O7WxaAgHrD36onbeUgEqkdA23
T6m47254SIPqAKOGVy3ZtbQOarxKIF+uRSN58dIXuDsZbioLuaPdlDYVmCdlOoX0M24fHVfv0it4
3v2JJsT7MmCVSPwKQdP+0k3JLQzOGxf9WeX3bQFeMlnbD16tQ4EXKbluMPfHkCLdmpK8Qtf4osiG
+NAjsLC+iOYS5U5+OM1h1/g6rwHphrMzAoQnRaq5K9EzIA6DI6YdQhwnEg+rE+YJG00Pf6yf9S3l
aTQFRC3oTV664ZynImyX/LsoEh1LnIQdrm8EXmPDLMieZtmcFC5Z6KveLxWhvYkjRQwDb1CeS5WY
RfgetW242AZvtrS/3HmF99JA1AKlL+BjFr+3QI8fTvmi6ymxCDOdlSqyyCmUL8D7yipgro+2mC/K
VML6QFrfL+iZuPqjScBmOt5qgguy0rxn15AgVM8AeGeGO9rRHomqKepbHARBOjn83z2vjIFSbhsQ
d/OJMpHmDxvfJiRuMVN7viSZA77tci7vi0pzH8wCAbLSjijPDCEqMjLbxrOM2M4aMsT1yBQP100H
8GdWb70ThlCfSw57Qj55cpe1imPG3n43yGs3OhmDRNm/pKn/OxijzYQk/M8cDySvTS4ipDXeDhQq
UBqhUuwxuWLfB1CLMHmyjLTtvu1wPhpB/4FtMe2ypCqmJclsm1isY6D2eL1iJmYjd9lAf7C3kpnR
rqiyE9GeBvhZ3551Mu8tcWTLzibLLQHVevjaRZW7TQ+zV8OC4Feot+ZH10dP1dyqglzwiQD2+rud
UhtZqdLx0aRdhFa/khnZTrdHWayrxJs+YcILHcawUhc+Nqjx93waWSREwzRofk4nqcp3YjeLDRjP
i4/9zEyiAiIAbDRlrHjOwzlKzVVs6fqzXAZhZEqZEjqbFQPuTfwqvPxIPyPqeAFx4KZuOBsqFEg2
8YGSrY7M2+KUQrMOidCG3/SoQNtUkp9okJLiFWmbJtCTLcH3abnVfv4fvvpY1BlO7PgT6Vq+AgyZ
FCNuDv+JfoWUMejnjNJaqs0u+hwhy6e8OVsyzQHOUZZ7LuJ79G5DPAEThDm2j4S0moQwZuMr85RF
NUl8yroxHmb4o3ovNqkkH+XROSbTqLpGy+ogZq8jQnBNIAnwFSAHHxIj5cPCUKC+ea2JLaYnzrBg
/WLb+N7Bn4XWQEcATPONB5USpsu2QGzg5yaBFkZDmMuKR/X+R0Q+ipYb/YsxjxoOXCvnbm2o4BxA
sQpmhYPk+yPMYYHXS7JoVteJ8kLCsGy8lrCho4XA4pJqpZZX+fyhTfZ3lGOmIIzgt75bO3qIPMIO
BAXTxO2oHrtt6Dd0dbN5f5jvSB/ms4pwV0UdINsDe3EMLZHMrR8Whx5/F/0cw2i8RNQsP2YjFCer
vzhbDHer/O0yK69V5dm7wEk54l5VB8FPdW49c461p0UVGvM1tVAg1xaUVoOkRrr7C6n8v8GHNGNP
mFDXmqPbN63RAn4qeCWLGhIXJ8G7RtATek3Xf3bph2MfDKXFTtRFUfAbBaWHhVEFj077Ux32jLyB
j9hqa0nSuKHRAQoGcVlEN2C9vHLHrDppmBbHcRrh2A40IfDR1tm4KbZ0MLZepQyhxPHMmmuC1G0G
jLj1WHK3yVMYTXzxE15rzPUFi291S78sHbVeFwCtVANPyuia5c0fqhp+yBqJubapyqo4ww+LA7zs
2424idmzTVlhuLNROFAak/9ilkeFMGBOK2e0KN0I/44mhReUnKIv+HxEIPqRMCEZv1dwEQRxkmLe
T789wYwa9iOctKqn/joFctz/tW7OxDJTqSbff2VTZ+dP8Tu7VVeltKl/zp36Pxp1lfH3xjYI32zY
LtUEdPt02Mzd5CE4MGxD6e2B/pirDBB8R0gKIlA/zFvPepxSTkWwBS9zWyxsVLkKDb7Kfxi/0Nk9
n2tHcbq+hpyBKDFRCGYCI1IDeErnazsFSWvGTCnU/nr0eBZrZdURg1ZqP5O4HF1JgdrIZ1jVfOqT
4XVu4coEtZx9eNL13yeggZCQqXe2l8m3kqkWuJ/9ZQ8b9aWk5AlnZwYQsuJgF2I9J4UyTEcBMVD+
WnYpAvhSn2fWq4zXQRs6IoCoSXG6Oc26FW4JDZJVjQihfyXuYCWrjInFr20FnWwfLMmwN/BPHkIJ
JaRTWqJWWEouedzUbYETP93k/SJTes6Z2ZG8SXgHHKHGkqH7J3IUuchjWGouX/2tignU3GdhrSX6
KEnHHTXaNXp5+X+k2R9IOoFqE38Txe90sGOJX9M00/KHOKBJtW0eTj7jSTRR2nE6oYLLAIrG5g79
0Hg9AVUlnH3W0VOOJa76BEBqjSmcgMZ8bP17F4mZYFaCkqGmeK/6yCFBQQv8xzrT2P7tuJqrvsRj
gYjAJE/21wFJNw1SMwcggz08a8T90f5VNQ9H5TJM97gUTL2QNn8c0noqy1E7VpVEOZSr52TKiM47
vS4ZtRs+1qxg7xfZcy6boehhqHENFRnmBO70cxICEroR21bVhwnDJmt99xGcwIambzFVZmZvGjce
p2nQjadsQgxoAvJ2usyI7DbwDWwNbV6dvoHe1ruo6+wgmtCNPCqyzJmzJkNKhV92Tem7sauzWUce
9xCt3KFQHx2IwTdUHqQ1pMLKAHwo/G8e6edxDALJMkBdtNPXShpzXtcJA56603Me7YlbaAuipmsN
1ZpU8E6nb8hlS69CT9h0BgdivBIHTK7NlfsITpQQNpW1xq6zD8WISaSnB//iLd+07LE7dJ4WFUUk
uJkiBYnk1WG0krArsBBCM/ZIlfc5f9/X2JrFY0CczATUWmdbF2GQtxSjyItSyn4JV6MlCAKEdtF+
GC8i1goRwmYOeLI4lEoaYJX0lSG6XUkhvhsP3A3XBDW/ebqc6xM35QwWqMatwpy7JvB0Z3yioJAW
lYp/8OP1sz9GNGOShiLdy77QyHmTpH6bTOwVvrvbdyjE5r7IdvErl/1CMwwYwLhcdhQHnL+SwzNU
uc+IRXs+lMFzgGbK7MzDwNIHqC5pxXuxm+NhY9dH17SNT4pbt5FOCnyxM5uNsiKQFhvpZzJeVg5e
8kCMRw7ACLmpf+yx2i0O8RsPYbEoCWreQLuFfwy9akIXzgqfsgfv+0pYcTkDA9HyLUY7SuH0YGGi
yxjZrdNJ1yWYPyVVqsZHSa3O2Re+Bl4TVFAD33ysLCW3NFwL76cL5zsMLjgam+M6asClcm8dHOuE
K9i9wR+m2MAO7Cw+dUNRLI/wFHD/wZLb/InIrXaWPSMVN8+RRBHNw6EkapNtROObtU9OsXzD7uFo
l7z7Hwhel1muaOKxAXF8tNdymCNAlbrFSuF955weUyBqwaVjSDFh5jaGkqCcg0zjKFHZ4XJa95fD
Cuc2Shl93Qx1LjeJ33QLZUnSUk05JCBVXq05z6sFomzDKVcVPqVAccU6wiBN/RDtK3jzc9CMAeCk
aqkQDsWErV30Ko25T5QqhfOCKmEV4v/w1eQrrnpFhRHOVPwVQmi8dVekn5fc+Wjvk9J2i6kA3F9r
skvvSxaXq8pUOwGfQYtQR3RVG1lFWLyYIq0wnYZTdSqgE3YKgxkcS3HFRpFuxYsvnqghQLEWOE/2
jnnUcKf+40C20yMsp64DSUkG1FIoUsVkvFeeIYWNTlfXjR95S2unRAfJgUHzmPGA7u218Ray2fbL
C5TwyzxlqIJMXyPna62IhxGxNUI8E3VtNPkNGe5zysVSlEqpDxpsv+jLfn+Eq5q69RYMDowJUgrW
EHtCw7dxvWWKZLlOpSiDoa/Pbf7Fy8i7Wn3+COF0sxA2nLMR9fgFVgPf+bZEwddRSWqfN+ZJBCIl
hDmC5hMwNL2PA/iFapUZNrlYm7Nz41FgkCQkduQL+OG0weyQHh0rICIgHJNvspb/zq2GPDfHL3sW
p2vH5L0UANWI7/a3khH8HX1tEuRMIgWEpEpRq5ozsySn6fcDU6WhTKyFIDhNH3UQX54sOu/XI7Uj
1BMa7JZgpnxibLkrgRRsqWUQernzWvxSnkDPSwYayP0Mgqvu8witJaoXs6WCIRJ+DUARJsZc32lw
c69lgBkTOqzWLXujaz9EKLK1gOjbA0CdcrCc9EDhvprt5FwrVxOz43KB0+HNbuFMMSjwHk9qbmQz
86zjer72cgAinjCiUSxT+YcPUPH8tVzuwscUZYLDRh+4umrJpCGxZPTwg8A0oiitpuG61DBf8ofK
lQIk8zjHxmc1Atp3byi9Qis0N9yXxuDZvO6W1/N7l2CrB3ZeqzpUS5THFYZFdz62ODQSICLBJzl3
cKish5n5R+42+PpUtsZMMxNI4QpbroieSZCZ422juIidOFdDf44B9eOI+KueUSkHEKZDPXiq30RQ
b3iFDriqUzwLawZZ3f9DmKc2Zbmm5UqNN5imeY4SNvZ9iQdbNsoHr2A0m1Lx7zR1c8gxQVm38kWR
xjUlvO1RBmwjY2TTKxb8u3Qrw0PLZqKJyo7dnpNayGF3RnXXyH44akd4O7JW9CxuC/0ZgDSNB5Y0
XY8HJ74+VTa+9kUkMfkGgq3z5Z911p9iO9laRbx6M+9d7j28cyrB5hk0xrYpHlNF9Sw2ellcFVPn
1taOcl7VsciuLHQil3g+Is67V6VyxjE+AYxW3v4WsFGN+zrau2VMwDcSIKSfId8wZ5pgkVf2gaEm
WBckArvfujl81+FQO589s4b0JLY9DTgwyCfvBMSPl0CkuhxHD66CjKaqOuqG3RR058lSquK+NN8u
cET4BeL4MQoLrHcb+WbMT5ikytRR9IPSasFnYcMQuJj0VDpJ2yPGOhnOg8qXCpIWBZngNj/jMEZG
VU4PpowcPzOekUtajScZclATtM4LyFrm9f9QMlOQOJSloH0aYV04SVZPPseovTBSZgn7oh5Di+L0
rBzGOy0uOOArr/wBtlsWM5xqR3t9jdp5Iqyc12o2M8KMRHunX3Ik8lLJ5sr8Zk89K0/nS/q3SZoa
DPGrzT4nJ8ZfmziU0hyHK66uW9gBLZYP/F29eOnAkrNlg59gcbaZuGdsjuNHO7EtfVF1G/+qzJFq
J+DU7jLhEmlbjGrOn2mo9/n+RLrN1tAYhpyJsUvtNlwRYpU+E1XWSoAiWujSHZwqyo7Z+pzLvFbK
DKa1Zmp74S6rS7pX1zad/PgNLqfISimdJ25dJ/keVoZSSN43QhrafF4MZsc9mWt2WRh7/KUr2U1U
HOQMSJ8HvvYSm0e1I2Q647xdHzXwmGXTtmpzFfwjDGrtTYqq7ZMgwHPMaX8uLQtcmNm25FtZadZn
L3pgSNLOI6A5o8PH/S0q/xmlSNjdHlZnXXMgJ9Pce8w45uRuX9zy7Qt+yJS79OpeLB4Iq1pkVTqq
A78Do56FSlse3vgZXzprrKtGn5XrMkqixGRopi5cdMu4vMMCme0OIWn3Is5hSSge4nILeemU5hJt
Iije/BzOvUOTfP/DnUzuvSlWO/o78wAOSffJZZWLNMYD3XahzZOlD8iyszqDL3AntP75uenRlouD
z2BAQKUs5iRdaIcfryStZINWAPL8m9R7f2Rm04X4EbuL0Kx1D34OOx2h7HhVviqSyrbv00ZURR5a
ctOMm0g4/K6nHzSmOqJxAsckjjBst7kM2IEofIXT7PH5JPSTNDyIfYZA05Sg4zWQDv3ZAX5IroQ/
sw3G0zg7zWG0KGjDNlKEjga0F9KPSXciuZL6dPqvvG+KjZeQRtxxcHHRAt9J39XxxQDFh2c6Pak/
UxeYqNAeRJet9QYXohqxdjymhcDLDfxa70IG62WyRQE13bj1Al5e/WRF/XA/geb8KwynbbiQZA1V
pmkbQ37tJarCsB6X8E8NTIgimzZfYBhrzUTOp+7VQikUyFRD+UDKoG8cNhr2WwqfvZoiY3UCXhuR
WQUdbr6ocq9eJ848sj0dAPANdEp2vsNcZEZI1JtshDXzO/WFTbUu9iebYHq7Re4Gp4f0X9BWSoJv
fMVG4dC0DEk2ioxeuoWikO/kmgMXnGWuJC9r46RZVuo7mua4Jb7QLL+A7fiPcSpFYgHhveIKohML
Z8Zdpi9vr/U1XsOLWTjz/r1K5zhZFZzTZC0gz2f/HSw4j+G/a8isPDzLw2mtUM7l63pOKPx2f+Tu
5RVR5FdAeWeXw0wYfLoyj7J0qYauvWIedlrxy0XwD+NApq7oSgpYfxGqcSprNJnY0X8Hgv12nHBH
z4BnHI9KBmXfCwPYSp+FJoDLw2LBNuMXggc2E0nlbCpAenQpG+Q7YWo3vZEfvsBMkq1hOP6DWsAE
dH7H6QSm/e/ELU3mKSDCPaqk/LuLCo+AAajp7iPWndR5jlPniLuSDUJCV5xi3izdFcLnndYVz/gU
nESdNqidr4pytzEeGnVT1yi6+SW6wIR6SwdYu9zGyWSvZS6egA1F4x2jir3ZGgAoc6fEzMg1PMxN
cpP6BoajRAjR8ExAuUc/t52SyTS+8DGGy931hS3yg9wut/b9FCVHRde6ZxjDmnLiJjwmd5Ym8tx2
cDHgcuuPj8+ScN6EATVDJ/n9PTRdT2xRC9YMsvrfrxyEqlHzxCo1sUrxNT6WmXJ2JcXcMfZivFqi
xoSVuI9A9OaWv6gzEzov9i62zx/VKUxPgwKqQd9QiX4o8zR+SJLSejsV+zo815iXYKjcxduYvzwZ
OUGfLn1rwdG1kNmRfGr33yYLEdO4HHz3cLll1+VxdUr6Yfz9LjP78X8N77+lDiB43blKFwdkfKFK
q0CO3sKm5wWp6Bi5a9qwJJEf3XJsbP6Wh0G3hmCvf2/iI058LxaDzqZTU+XpqVpjrRZMtOb2M8j5
4H+FbfpWnS/W7VBxbmQLI28cfVV0pg4a980Zr9r0zgAPyWh5WDbnel1+X6vBUMhFnYI6hyYnWahr
nsE8J4O7kfzlzXqNz7h7EvOhztkuhHXsQu/zYMJyCFQU/49AKBeUHhrwFTrAeaaTEiSDAdnMLwIY
SP+iSWVIyIS6Ypkuo9gEU9aeTBtmaywQog4Ipb63Sg/WmbV1p1ESEEfJTW0lhxW6+3qUgxW0NJay
lUacKBLkryhCTJnOipzAotXPMDxy7XWsqOZftMwPOrJTEnSK6J+uL2ZdVG5coCABkgke14MxW/CT
QtE+v5rGt0cq/RVPxUNSwNCYzDqPB1Y/tlWvo3YYMk6JQgUoZsogki/E7PKMaUf2KWsFDj0ENW9s
wO2HdKd1EL4noHkgZqsucXJhrEpfgWB/UTOM6lgxC9RNoYz6QsctlUW+p9LAJv5gERwveZ6wN+n3
lOcqdrf7fYkheDP6wVt5gSoz9Ytsy2OZ24JZ77Tr5w8PCgKm1i1js9aZt7frU6AJzu/UPYvlkNMB
44Pkj3wolNPoaNXJtXp++KtzzCpRI6Z0PYWds0iZtuFry2vASF3pJpT43FpO2DLnNo4d3H5opE6v
hHGdFxqLHU50dz/TGlftjFy9E8Xv5hTluDTgfCjVdVT9SfUEejkyuzeB2IleD3ZAq5syjCSmXNmD
YV6YFndxz0RC/jyXyg/OHI03I/b1ghO2QHogBEeetuGLyO3K5mETbwo9nqOUwcwRFFjo27e8Fc+j
nzNKzEysY2Et2s+JMyl7uvUwF+ZBeoafRPX/eRbIJz5qcklqd/wiX4GukOYlK+qEImXAVpC7AHBy
z4j6dNDqEAI07lQ0ga/sZ7mz61iM4njAKbUVMAhCDIBuF4BGmoLsPjv0sKGo3lHyKsJ7e9/+8PZw
Wr1Ib8oG1zH23f0fSVFTZa3gFHfy6H2/i0cwcgN67sRdBHrXQCTODDZOlPN5avVtkLYfTHcdTYb0
lJLq6M6+KnD/uBrf3XR2UTjn3Bbb/mE8Kao/UEs1XGDzTgmE1wsOE9BIbXlaF5u9UPV1feY3m4Z5
7Dv8A1vnMjuQBGdq4NLiu0Io070N2MvPGiGXku1QsG592EPykCaDNK0HPiIvm6wxMb3TQ51z6kih
MEeix2BRbtBNY+79ngnPXTNqXemGRNTM9pD4FdOjKAW2RumPBnhkSliJxQkBWrs0LjqiLM05NJ5z
7GpzhxzYEI/hRMxkjbgMkjwQ4SqZCBsMKE1a7eF6G4zY/FQAcUcdcwHSwzGE8yQQxWIeevI6Elqr
csBZh+B8O4CoT6Fij/azQ3bgAAMUUleFG6foY3HgvTwhYgdhQdb82on6ByM3ZB5a3EupZteS/Xnn
SImq5lLCkGOFslb6gzdP/R8NRs880RKkaBxDI5ASVEq2fCOq59tpdUMHXSRgEw+WhlyxvXcb/yF3
2aSfpGi7r3Hedp1MH2zED3Z1kHnvMgtAuYFoxs/pjwvxDzP528wmCq5NsEgAIzr0d+kg5OsRx33m
m9tbXqrelDYpXgLPNU3RjpXEjQSQAlaCacuPglZioQKqM/FxbuJgtjQotWfHbsRvMFmEk7bqJtdm
lOT1ZG9HiWu/6jgjm2hu9pU45X+L4E+HFcr1qA0bGR64IwnkuiwxM8v+WbhBlpGTQTEqO9J5/WUp
mZ7VsA9gTL071QrODHGDt9LTDA1/WKyGEc24e7ayzx+P7Ss3qmnC2t+KWgEHEQQnS2M+he9dkS/N
eIVx5+uKorwdF/PcmIJJ6aUoVyXFMybgC5qqPkZ/Qy6+SI1gJ/hK//3kJMJQtl6VPqy1Zd9x9iZW
ybTzDiU4R0GpiY5z5pE82sR2idYRP/7xdSzoJ/AVubvRfSjZRlK/Gfnp8oty9xGTr+9hfxQomztR
iozFPrbruuc7ZC/OCd0VhSJK35sk5gYnzmRtiw7aDG3wcWX5fj7FOI6U6pitnYHQL4oTwPZN41AQ
B/1NErVvLlL0bvSF/Gn3mDr3WfPK/Hc/wx1iXvJiSVeZyhbJy1uBZ/F+VdzvH3d0Og0cmRWmMPII
NSojwlWAEpiIDrdnJx561yrYf3iZZYfTRR6VxTyTVI8H5Z6skNLLI1VIsiGDfVBEkCJ8J4i3dUue
G52mtVV/Nuz6zW2A7VsLhoVzrLYepPMJGWnAF8OiNA+nNkSbxaEzsv4ddTWch3pUc6R+3idJtLvt
KpRg+GwqDw+zvSjTJr0LTI3GwrTbRfm/uBEX18CEYEfCQeXSYz+f3sKpT7kvYCXYDfRzv7xMAhis
20cY1UprlgnS8IhHEzXo98fySpsfeIZmZqZjoXb5/GsB/x0Szixo3rehcsYiiTgXe8Kvnxd27uWp
ATuLtqnz48VQ9pFmfMGgRkn4tEbD2xJrAWbteSfpQkaUVQiWGdP/I6qnwYEuv17Bpqn7UJj32UkR
HDbyj3SZOUTGbhWE/JdOyyo6adnBSogsWx+RjGfYfrRyQA3Di1sT8YogOJSWTLa/xz4XW+62K/uL
OQhd7COjq2sdxlNhvYm/48iuyjC5eGW5TWMhJtJGZSOQSTfNVrGJ886KPjUuvjanK50d+6c2jl+b
pb4XVCeCEjIbZn3LUC9eQUh+J4YL4ufbX0piKsOGdewlNL8F8ci34xfBOca95V+3PzEHoPKhinN3
2mehXwV8hjnEJhootd/61BP0LXROEjud59p8fpCjc/Pk2AllsVvA8jGG4PoqnuQng8+xhAsWmjKj
QJrqM2fCUuUukjQVB+7b4gex5gl4yjzUUllDf/dTcUS/bEieYIUiIskktYrIF4YXgjYCz+qTe1GT
uQ2NxIuPOpRpyV79GRLcs0VR3dwtKSP1H3i4aT3ueevO++d5kOFFhTnh+wRFT1APPbamroSjAdOM
yjhhu6Hf4lNCQPBgcfLUqhuLB3PXGdLyv6koXPkdfrPsOHg5xjSAHuI2lmohY2Vr0C/+ahRLs05Z
d13r8h/00yOQtFJyWkjyzZV6uPnNoWBT6VEMqKOV7wt4g/kBEWbT+x/npSN+e1YAXZsvsa3zTukj
9dT9jiv/bzu3IHYI6nv1MB6zX5dYbUWsoWGu94zuVFzZsJOpLOlqbdkFLoLZX3mHT+Ud5UkRcTvX
n6g9KW0knPm6H151Ph3Wq/nVZKyjM/SMNnLNREQG0gNGzib4e2jRuwaozQpulH7Ao8He0z8EboOW
LifhVlo7vdGYJ0rHoGWtjO3TmSvUIEF1lgxQewWcVQAKxxcu1/NTOpOpNpCV3s2Csbz5shfqZkEO
dTJsCTgLHoBNRCuVcx2+VgFaaFJh4TBtMRMpUebAQPZNEkaeLQVRGXChFt/q/kmGbgh6FAm3P8EL
K0Qggap/gHRCzimtIOfjEMaxB99z7KBrJqRUiY5csE7n6nCVWvPkw3CpXkcPcELMIVOmpe5Nlg4N
Ky/YLgWfyqPwz12mWlVxMtQAK/Ms6DBbcNwFtQRran7Dn/x0PfdTgvBnpCEPdvbmYgDY8dYvK/x7
yx/WXN0aR75hB+AwjaPXJNILjNUhq7PJF8Ca3V5k4qPh71MERKeV/PBDskZv8auCRony+RvWzNqA
W6Yw7/P4as63MT8d6d5BiLRAEhTISyT+Bvn9dQc7C/UtqQdTdp4Qsq19kpGcNuA1AWtqofq9gXed
6nQe8aUDhZWsZKxg7JHGXL7bgCyr9CDb0MFvDVL6cu9TEwgTOPMmDZfkLyjZtjMxu71QjVy01whO
SrU0kIEflevXNbiav9FcDO4mIT9Id6DGOWPDp2S0Pc04CHDNhcYi8ggoBhKghZGssjrSxbp4br+F
r+wb8ffhmp6XXPZ6bxG9Ybu3nVyjmRjucXjHyvUApe1asoXm34gok2gwylhY1Az2z6+x1M+YPFpx
dDM70Xy21NaJVPpaQGos9A4hl9LWRzhoO5I2B53FJXvMXjUShJjBSl/VhfXTwdclRFe88nM4jpVD
eRh8a2OMnhfO6RnmTn6grBH92/T2ut1AmwUIKCyrQooOneCTNr9s9IiqR2olF+Y1Fmti/Ap2grWh
B3b/lcDelbgDNLinzemUM4vsrrQQUmjbHgUoryTb3hr0oAuLXAGuX6zJhBiO7l9AkpVG+DWxL5zM
vDnP4LfPzZO8MBcrk3vk+RxjX1hsqwVX7WZIYgoezxR9eoKvadW3zTg6HsaFTv4oo3vLGNhxkn47
tJVzQ7G0o/z8+JjiPjkTf9yc+ryklpMW8Dv6spL9RJJ+FzCN8ySZuqf4IJlC5sk0ViM3qT9v265t
FmAEk/YrZ1Wq6PK5QVBZgYlXZNL6aHO+iX+lFGgyfBENa0nWvEtyTswdb5bDySNKZBuQ5ov7j/E7
YVnM6Hd61c5K+UgHV5d+0HnmdYPZuwGQgkVceXdSXyf5hFCMYkdMasGVkGPaXgmSkxAEkPF/S3pi
BRXnZeOvmJIX0MGm8xoVcOJib0ELILW27NSN+0zheK1v/cDvzm5EDKu7zZYKRsaM3L9Yd+mJtsRI
rS9GF1mCqqi6etDdEpyICz8p4fuX9VMNJIRY0Oy23ahMI5FLsDKKhNcOjG7wV9u/NCCxEUT31nc5
mg8mCdo+ugaihOxV8DD1RKXkCztdr5OqjrdyhWFPa4O17IJ7kB2riJInZN5hlBAwKleGCkDjb5Jh
L8Pbyt+fhZbKguk10lugbe5IOoV6tNbwLsm0e0jW9uFdDnF/Sq8t+GDZu+8traMXxeUsvxW4a6LU
sknNpM7eTCUmpqkjDJxa+ROWEOH2bXBktGn/Pp3Wls8LWqZwEeyWpXVn9uYsI8iRpcd7OxZqBzrM
nk1Yo3rtPkTyX/gTBgLThy2T0Gp28rbMg0WUV54wjvPGHNmqt8Jg4ftv2fXmi9EnfK52plVU70i0
PqTZMIws9+p3ixG/JcJiHlpzakSJUqJ94TLAcMZfpfDqEf/5YN2xJfae31uVhKaaY1i8sjFSsb1b
RU6LKOn4ExBiu++Xwv9j7oriftC1gxXGL5Wq3LGbmExGySYWFw3DakHiv2lG01Il+jXGbX9pKNsN
Onoacv370BDHiOB66JjSlLlNvsqRzrBXGVXZbZzmp8uynTRf/R82Whu5Pj49iqm/TK9K8r9f6uK4
ioQ9E4ACwWJFCSaEiFCfyY3vlZlWBOJSg6exZ8T4oCilsbwiskFv2x0hCbObc2Wdo5eroE2dVxx6
HRZSqiFMAyztwzKea1olaW2ak2r/40QhRugjdNxTILfOrh6IShzroIVxha6vGYsWynRL1ddXZe0M
lz7zJRzU/GswbpXGIhyl66qnT3NgClU+pxSaxWbc9KY29FJAMOSFW1KQlFhOOuqBAppcCldxsbRq
EImHPaf3r2l/Iecjh47vNrkjQwOdciivDgNZPfZ9AJXwHSYoruNsADYQ4izTBR2hTzKVTsQg1JCI
quj8LU8X5WTxiCde/zQa8dNl06t94HXvqTM+HuOBJSNV/zyIUUkD6OEkTd1f3JCAcx8OEeGxBzHY
OrCTYjbCaWYL5UBheI2y2vy3qy24kOQITATfsdq05uPlibmQ2T/pPNULP+C4PEFzkg24HnN3KXbV
wTk5xgj3rgjSNyxX4Ip+WeyTaT3k8RbIwG9AGZ2T4X8qbF0/DdMrYXwXxJzTVvKoxZhWhJAU6g/2
gsewFlt704JqXwKVsUg06sWkXXLeSfvz2sCT+Wsl850GOSelyKcsOWGcQzE+4uZrUyFxKgWn5PEY
MNdrz7W0GhSgbdC1OyEzySNeVsuDr2dMTTecImOqTPsiQavpFdSCY+2a02Qcq7EI6clXESXG9fq9
BdDRG4JQE3bqjoFyO9W2Xm0Z48r5kXLBxl5rFamkjZBqzsu/dI3M7RFMFEALhRUNrTSEz4KFYG85
CF3vto0k4ZNxqYHq3MjurJY0vUcG6zCRyRQ/sH5jUQHEvCkIqovQlGBVvQ8lprZmV07kbt1nfSTJ
DTXgGLgvkKamYN8tT31K/rAydCzmgXpVGXI5eCI4XR2hwAdmmaIDd10jGadVr1a6eiDepGhw9TMU
DH1jZJNZ3HpBkv6eAGsP+8Ff+GytzOKJBNUKIncEX76STjmO0p2REc5dSfUjNNRuR2jrtl4WKB82
yWaOopX8q74EunVqv4ImpFZ0eTaHf/GW0ir8thTrQBIEzYcIxYeSlUvkvARBt6LwKb2XgLWM1AMj
iPDYojVNWm0T+f5nmwmvNTdTgZRE7SDlXkFtuZfXEguLri+AiWEKnoS2ypCdA7pJH3PZ5v08vlZn
20EBTUMePxyM5H3QBhyYW4Zk4Wi38WKGCfRygJJIunUZbei3I/UIm8i7IYLvwQSW/CraSulv1Ol3
wILRm+uCGRnu/Mx1Bya2SCTolV7jcN9nLdM2M5HiFlVPDRw0gj19ooA/LgHvsOxrW4DlulN26mWR
LEgvCHhhvMLfm8TIkXCHLBDpoo5Si/Wgawfzh8oUibR8E/Ly0W9YPHS81+zOXS1xefFIOu++R/FI
6DLlB7fop2AKd/RKZTPvA9WtpjSOleXJZ6K0Qcxya/Hu+AE0vNkIxC/j6QLsGkpNaHPFfK9VZqW2
PIonlucMNJwF/621irss612ZGnHThhmUvO0qyQeg/1JNqpubOXQTAwYTY2dNpzTt8QWCsJMN7GbN
l8mNAEmVIPMSfBy4DPiKVv4rZmIV2Qmzbkcw0lhXYakZ5l+zxjHYeC8I0U+0UpF7yOCqebvXrehD
WGs5H/f6uIyFsEnyv0L41OGSczYXU+3nSl46M7SOG+ScAk9OBVJ/o31t24yRMmKUJQltdvIeZGgS
vpOwwcH9JNsQNQaFS2zlnGj2bBbz4chhGLYtCc9Tn5faEEOaLbxcBghTknSN9FeNqywUaiSlaV51
I6OI3qiIb9WWVZZdY6ob+xAWAUkBCqE2YZCf/fTr1VHYevPF/O1H7IJnE+Vquek4xSoAWfB307IS
+2wecfIT+an8IGdzowsCbCYUAO8qwNYQq8X33SSm4LvuC958t/hbfnxa2t7XkH2J8kSSCsYFRd11
NCa8LT1rUmfLxS1gkcu9+kFAEqpetSA6NU+Ohxm6tajgxV/54l/QzUJtDyzNDgGxZHH91WEGWC3p
fqgVZ720ywnx/xw54qA+tetu3edh4dmCIoKdrIHu4O47SyXtprH8Ib9PtAepRgv21zzoox3i8a7i
+q2PF/OnjV9FBbOQrP4M+KOAlBFjNUp43+bwBwhnefhiG24qsfnwFGJw9Jt6GTpaJcWstdugUERE
wvnTivk6UkNHukpEW720NhCGxpmbNgrB6FXc5S4KQpjSRPi0Uf0PZ3NeYN/413VNod23FG2Lhsxf
3HBMm9+qQhjHrklCRUzKAxg2JnfDRpPMDCzrzN+gqAb3kIAhXbZ14//IPcu7e609U5CqfqrIyRZF
ee1DWBisOIOyRVq0ysFLjCPJwBVgcFXlOvNxMRgXoZnNmNWXNYi+HgkBVBTZ2mChLiu1daBYycPo
5ajYMCsgo3fLUciERfelv0qwgBQbXBHyXaoRyfL1TgP/rP9pcgIgr6gu9Eh/PmSMnxBkxjscteyW
8gAsZeKLF0ZSMJsyLtXZrXsc9c5d5yn6LF3x5z1msqsBtMI82W5P2mHKzrE9asckyAICFCJJIoqz
AWkDT6au94ZLYVALW4MvGe/LlUreONFr+aWG7SwUtfVprqgE+HpX6Yj3QX0BhFvbaB3aZ4HNmlxf
wIsC99+9O/Rmr3MqjTUttf/8sNavi0epxTmlAq4vG1OzoW1A9me6bC1cdz8jgrJdjh3Qenuq/Qfe
PA499TmgEi7cBvmrDDcf2hpclespvcusKGO8yXpB+yRHGxjRv4eRhJW3BIgW3wt/Nd2uokE/wvlm
Di8MDbrsphoHat3Qit/RqQiDULETZa5T/YzlWLSdsYKayv7fJ/9/bC0jnlO8vsjKaG12eAxoTjTo
l2nXEbrHjj1D1qCvm8ieVOHsTZAwX13LBMuZH6M10kCkm2+Ed4tJDfOLvZ3XGW8iwTaFSF+ueX/T
mQ03BGaCt9phDPZWbTLbh05yZlqD8mxgBZHZ54VDVEmz7xcQU+o1o3w7A2wzDXvEoOr9sIFCwmFP
bO8ezKFDO677TsOo1L4NJlnplJypFusqYITEy7qIhZdzbMjC+Ht71nBe/odZlHNSpOirptSIPiyG
vAhgESyovcvC/ZEaX7Ua9MRFcRjsC/+ilq0t/2ao5OS5u/m/8AwaCgK7urAKi+hu+GZMQMxKosLE
kEWYFCi3IuB2zkl2MtSvZGlMJU4g4ucsGNCXg15a3KObdP49TXq/EYSPKJpUYgdT3Ocx6aGZb9XW
eFSr/iydQaeQ/Jb6xMq62NTtr1rhWExVcy8KkgFqoA6lWxmZzrtihhAFSdeZq/Lx+m7oujbB+/dr
1hO/VfNumFsPvrJliEG0tYe8cOeUCKN3Aw9GmqIsPUBusCKqBoS95LObK+CSHfdOXFWP+GhqKFUW
a8mjqwuqE9cZYJOQU6g+UNgzE7YQNACrZMil3yQC0vQOQAkk/7keAnolLxjiU8duqr9EdGAwuThe
Z3spZ9ldNVZBVEnWW3A6+RiyqXn4TG98MhBprZFoYDe935ou+RtAJjg3CHGB/PMh32ASzBJoc2fw
qbVu1vGUpWGiVrlmdCkQ6c/nkIWU/+c9Hd1QZ+mZ+Qk32UsFZGWM6BbE4A3qFE/G29rFT9bg5rAC
ueqVKesINC66FRbn/B7mThuZ+dC9c2Y4HQZU7p3JYfMASWWsPSTmrQ8qZ25uCXolqA4wNB/AnEpn
E4kuyPWRBSNDXLL0pVqhWR/BQqzBje157RyISUHpw8ilO+g5YFHD5GkLV5KNJJLky6DmzhnwYc+x
juugoMRy7lwusXP4wMcM3fUO9QtQkDzujQEs7hvdgvUP/z3Xwy4rIeUWsFMC3/4cdMDoEWp9XilI
CLrCMQRmwz736Xkdsx/vvMyRsXNtVWcls04b2RMBwDiBEaVsJX9GY3UXEzO0S8TsldosyNqjNHpB
p9oqrYV5BxSknW9lQYpkK+KRtEQ8atDiFE1OgmeH7P0Ixjjd1LI7kEP9givTjrF8jvWXmUMLBOLp
bnv2zkOlg35z8z2sNI7rfUv222MSnHdw3B0jdaDO4S2aKha+AXCZMadiOu8O1BsE0BWm1Op9olcF
Caoxa4UuG5mBFWsSR4x/lMrM1+We57VHiXOx9AGAGipFCICfvloZSVywv3yx2K2fbH/j6c+/1+1/
4uhQotoFQcCQ384IqhBaO1ALJdZR6r7gKo9yJMh7gmoKboSNQ0jW1qT8Z3f5aFUw+/F7P/zBAvgt
XN2ItT5XE9x090D2nnXP/6DzpW1920uGyRXsQBtCNwwmtCoNLFWEP8wIQzYKu1wAfa9amM9R5WWU
DAWg3rLTpS6Ut14zIFvLaBPw+o9JVvFWCia1DHlgGOhlP8NeoG3kHWHKeMo3OE2cq12adbvDZkvr
m20US9lcbjz7DnvYlLPpyvrskXNaSiuTJ4oIbpI0G6oorxtpxLnU2mGWBcVOt4x9FpupDbzqXEXk
u1vhO+IWawVX0bDNJl3y3HhwDkWrc13Rj1tCOjip+x7IxWz8ibm2/eBfil8oKACDPyxSJXsgpRqa
SDK+SeFPm0QRWd4WhM55gdy5EU54j5VNFgpkmRyg47nzk7nCRIjsX5ej9kZMmYCL1+lo7J3NGpxf
F2xNSdIEKP8VD3JJmbaoAmtZrzmTtCstISdAvKS8FGRUZHUp2CvG1qBrkGTWYHOaeLnmCdYkld0F
IFb/1eVMdNX1EhRFRAHoAXzDKYhf+UcGLQPX82xMOgGNIyXJiTyRMTCIegO1M9MEztd+vQ9G2t9k
ktHnxuPutAeS8Wep18HGT4YNeW3JFetZ0tPMzVf8R0sIkEF2l3y6CigJOvpgYKkeej4JLu0Sk5Wt
208z5dHUyvnU73b6vDFP4e43VJmFN/xdyrMGgPC9pph3rXV0h16iBY9wdmslHenP54Dx6PO9Y8n1
0fp9xPWKiSBENLvBh8DofzGwAXYN6NmXnvJv8ptiUgh17sDnMBweA6Sv5jncvFnSqKbVOcX3fIUh
s3NEoPEzqrkq9qS2iLVdAuMYVHgb7Ymjbo2hHB2TayrWaidxaeywO9IdS8cvqG+yNRFdrl9B8iyb
sIGNcJXIFRguxotR2FDavZq5/YyK2BQwj8v3Es54KcPz+dVIBm1tKzegegLD1+9ifcxOP8k/Cw8e
kWj6EN73qHE49vfHqklk6lFI0wELlaQfGVXmf4SbNb0LjLLK2H5Z8Xw14JT2uQJjk9l8a3ynb20Z
bkMIvZQxQmc9Mz+Up6DAuW66ObzbJh+4YGSQaEYUNRneFVFm8IK+KerfdeDHGmDy6vI7wMPf8q7K
JxB2PX/bA7bm0lSw3LZVrpxm/jQTtMGgHc2jpkhvRK/8HglEJ5RuzHDElqHljR1x3K1dAhDGI/OE
PiqMGMUm3zEe/n4uZNr65xc1cnwawKTf2YZNsoT+BKZ21ojnX0LrvOsdAviT9WLgDCeClryfrarr
SJwR+9HREhnDlmE+WxAqC2avHkAyUjrRQdO8oMV8Ob7s8fj4FqcVIMh7jAGj/Y98/2aeQVa6MhkX
35YN2ZCRUGfaKTYRIU6C0QTyplfQRX0gcZmz01h0WK3fB3Nu6TcACibdmLMLeGLsLyzC2LSlsM+X
JQcXGDzbkvtS+aENsXGaycciDuOjROhn8upof/XVJEcS4IliOFW7E1gydIX3SHFliXXlLAIdA2hI
badIeqaeexyxrku55ZOeUHNOVST9eliwIdWFRlr+tNOc7/SGyUnajEU7nsohCZ4DtquhBsrPZjwP
b4wop65qA0z2TMgUzENaNOCIb+w/Tb4mbHaV8jtAT/iC/oOy4VkiQaCSUfhtD5th5MpnMb8GeiVn
4PHoiMw1KdPCqXrLFSurtJ+vheXEPYjsGA/pQMT5+34scUjeYxWBEQQfSNXWcChWyOeVOdA5GwrF
Zp3V5UJZwefjWN2ZGXXzSsN/GvfngMp3ZxOJ/dsJ8g/OpTclulsfmrPPSDbeHh7iWpqQnuLAigiU
EjD9VzfwZlpyVrXZYd2+J0TX3W8LSwLzjI7WUVhpMxVoDXFHY8IuVyl2ZacJg6RwR6Tl2i/UoAyL
K3YZ+KfK2KmkFZadjkWPWlJ39a55KTHy5rUc9o2rjVPRedv4wVBabaNRz0eqNUUqUZ7CunkAsKPF
Y8gUbOP4FOtcHcD4c1WZl6b084Yp5UMd5nRPk+3YiVD7xMIN75mstiBL2btg35QxaSzpc6G2DPsW
3FaIq1RRkt166K2xFMncs9InUHTHxV6Z04zwjnKiaKwt1gnGp568Ab6JOKZbHBqL6m1vSxu1lSCp
hLF8Iy+T9I/P5YuiFsvJsdB2DgF8A5lyGJIehO26jsnM0nDtspGvOj0reG1O8jL7EMe2xt6mi1nb
fK23pvIgse4xlSzn5a+Pd+94xWfBWS8adQMmBMfMBZNft+0KsKK1h4JYwQOUJL/1nC23Qg+1Txo9
CiedxPwt3ZcfokOKWxJo3GITJgV56ifjlfp6u2qGwkQw3pvz5rkvKqvz1qmY7Tmw4PgrhemSYS0L
Tyd3TtTW7IlvCfw6gRXURc+ow5OEctvNYoibWjTMiX+LDA8iAqiKnX+xW1tsS1EoRCGoZZYBlQne
jUq0DMwlzHUy9gKpt8yMgLUISVdrTKSHhhpFbhBvbmsLlwY2Wy4j4hNw+q3fsIaf0rTCIpiq4bnA
VrFfeXePsVHkIlFdkOgsNJ1yxzKI9AWQwj2q60Ueg7rBWExHaRH+gOuCXZouSDyH+3QCFb196BRi
TUZPKjdS4JelaPAYsCuszlbFq6yrIFl+V33U5uVw1KIfmRSxV64W9W+12Ze68veIKLbq5ZQ4fddj
/RYRJ/vwSnVPMY+A6WfZTiIia4QrYGpyUoM6NwpRzNc4T9lriHfzPHAr6WlAjSEvtbfgJz/VQ68R
aDo+7irj3GJORVqTnJmg60QjKnqYVc0tapWHA/ktYRd9JcwCzUXeh+z0lgWwlYYV691BVBj8Pzn3
a97GePVpV1fbLzRVHMMFaim81kiincDoM6a4jhtQNGgIDZkq6mQsYMqJIZUvmSmyvd3wkdnqR0yT
Z0PRpoqEQWjklJcyO+bfpiwI8go4bMQO81fxbRFQbkTxc1+rdl8AmdbDoG6HDGKYEVkRo2+ayych
rOS+96Wz0xQz7iNAClC8J7pXKb4kQ8OWNERKlgcvI2y5NteY8U2oQiqaGkapPHFMYXpiSXHtKOau
qV/itztGZficUy9VAGkYJdE8Rvx5P2NpCrD/eLx+cvppp9mm8jDVuv2NL1ZiZsgPo8EsfS50qqFI
AcdkmhGY1WInHcl3RL+Fq1fhtS477S4XamtB3yWqWVa5kn1LOWHqrP0ratw11pE6WjP9CZJ5NF3Y
8w/vaNhZa9MzX8IzW768KdQJITuwu1PqpVIkwSf31+dOCgz9SEC3lEM8b+XShl6+72W/1tvo+zzf
aNDCv7q1RhHx2WQaXK2VUOVLdH2kGdxk9oiROAMovNE7mhdOA6yw2gNmcHBK08VLS+PCB9kKPTGl
Qj7JqcuN653nE9POQbwrHZNrlL3+qm6+wTxN3HBR6RGQzAugd1N5qvyMXr0dIGjnWHnYDTOH6Tm1
D3CLxfRx1WiEOE0IXt6EWz1BZnuxVBjcQRuxWdhhRW99h/oBI2XeK2q9QDf3mIy4slpynt7z/wTH
/yz/NIvp2BE0Eem23FWxRFe16nIfeNWkvcXSJmb3wVLB3JSNr0t6HY8WR9Q0LCTZm6zfRP2vjJy6
YgLrf1Hrqcmgj0rEPxnUvFDdXdK6f+5bZGUpHwdB5r8ilZeQpKpHc6+++ude2cb+1vTCKoMku0qt
qLRKWjPgEiWceB2jYRj/VWbgEl9P+/M5CrIugTS+UuJd6E5vRwZEHq2mHHhStM0alJiCdmH6n/cN
7yFcKFlkG/czpr/uPYQZACCY0sxsSqOoggZzKyUl+m7uBSl46D9dw3KsnKgHyO1IF2CDOIJo/8tI
QZ5AlY2Kne1CiV4Xi7+5h95BYkvzRlmDOEun/pnF03qy/X+2ArN9O7X5uX5+gcZAO9qehq+53poN
/k63/E8ndSPeaO6a8nNF+jsXcREHjiriZPh3WxU9ZjXAvFS0dz3VUb2Nr03wwwz874hh5eGzPFSL
g1eHdQXqw5dwCW/vkt/XjjIujii5Zo5rmWtdcELqObLsfpyzdR77QTkkLqYGrpWdJ8JTxwFTnIwF
e+/DE8EJl6940Ofm7Mv6ALovOtTe/8xRFVPwPEBnfZBDgVRsInADNftA6xFbkei+7PbKdk0NUK3A
GvB6Z+iYCwoQVMp87wyezYROyCMluenurvE4Okl/2ViKuVFQhfesHSHCFI/n33/EeumkXrqK9GUO
hHeNvP4VU5Vo8BMFGpY7KHRDGok4eJvONBmOWoN0ZSEHIETur5I2k5Wd44ZH1X/yU3R+frKdGQLx
f6LpY9ZkvjHdo4K/AV0ekW591ZG5PNtd7dE+09yeH7OeJsMdhUAIarol0B7+yQidlBXghh3qzGSk
Kl191IlDyVWiKEk6PfxfhTggqH+bZXkkSX3tcuby4pG7aEJhrW2AJWMJbguAwoJANaDJLYVkp0P2
jVKsiF2YTjT+67W1Y3qCVSqxt9hY7SV0QgYPYbmqYDvYhAnc/x4wRMchNAlUEmecDzsLl0bwFQqx
NFE/yHuSw6qczdBVDOEWxhfVUG126SeA7Rq+AvLgc50A6Wtntp1x1vvNSPayNHtH6S1AAwo9aRRA
hpEYjSNThb8VZKM0d+AZuh673EBsKv9OSLpxeW9QSeoI9+JCWG+pUb6xPxYpqT/f9MLZum0rMSxj
x80EEy/ymeYoFYAURCEUVwckZa8op9BD5hde2OUxk+JQ9ZeMJ86uKGa/GYjpd/HDepk7ZRUmsPFX
xk9QEuryUL+rar43JCSTLZij5FdZzSmgBaLCdJ3hqQM50bwGalxy0vYQDLp32rzl216RoWJ0X+v5
AwPLdQGrQesU8o9043bWeh8jtjP5I7VLjU63ujYDmwef8/WHV0U5hJVvUSZFYKJsJnQtyLa6AESg
kDujopi4HzGVSdjkFml2eiu6kpWnpJg8UENT+lIcpS3Zg/JydpQslGh+bB+r0iwYddP3ERmTAljF
fePlfyUl6CEYLodJ9b7WIZ1aGdYoZ0sKMPdW2708b0nm1/5RiUP8sSS+eCaifzG2UZ7j1AnXAnhB
e1OLK/K0+wIlC+5RnFHOT8XujPU0MLQS3WDSdgIzQG6F2VIje+5LgmcLCsnFOU/6Tc17Aj9SwilQ
qbWH3X1XAZ6nMpnuN4FtD2RkkznqyM/IKmkzZuyf38g+1Kaf9xPQ1JhH5pQqc5MHj9O/HYwhCfUJ
04dz8taoSn98a+fcn9tt1sKIJZe7l4fphx5zbaATp5o3Y1S+H1l2oa2k6W9CoR9m7hdz4/t9k1mM
5+Rl+kp2t+kwhSsBaOEAvIAeMpnqLn2gscXNTy2K9T+oaZLb5SzxlUOPqMyEuZo3Q8wLZUACIxj+
UHP1qOHtDZIUYkJd5r6myjyUBEDPgGYf9aUN9YPUOMKuAYLCNRdDJHH3NOQus2g9iJu83eSTECRA
qSKK/aLvViVodrgi/XGDgo6EzhxfM2Q2GAagrNou5xYWJKObY1XdLF/VqmJd/TkDv9SqAfKGGs+x
/gYpPsQdt5LhwXz2sNKNMF6oxX5kxK0W5feh9gFmesBb79KLHk9HOXIls9DSLQiMAilBqa4sE/n5
qhzEoMhi3NOOS00sbFpoLd77ud7lY+ZwFUeTcc30mk5XQxTEI6hD3eF3q9hZmTlnim8yjvioWBpQ
JHizM50pYR0mWT/iR+uh4pCRW1t9DcQeTvK5kmB1pw0w+tMQZP89fD9KGNCuKqtUZfBgt3vJG6Uq
ohhomD5ZyxRM5NmAgyL1wLspcEYx+NdTEs/xZ0QuZmBXMx9d3UQ5DOp1mg67m0r8r29dyoye/qiN
7QI4QfSz4EMr/S3f6IWQ1EZp2sWz36QsfcwXewUbnsRdogvIDmNMf8EHbu5Ym72p/wX+qkiYf6zg
jm918Sc6M8C4L2tyGdF7yfmUvfJXHVMLzLb5HrTlBIYfVgTs/c0BbvIDY5w4Nns0z8tAwOweQbYK
hWesm+Xvhe3KEWqpAzkVTzkv4+1Rjk4rGJqdeAuGnfI3HNbTLrIMAE5MCP673ymbBbMvQwqMCIWA
5Qgjnkwjs7M9BVhTGZRnSFUltpbS5anm0UZ5eoomWM7foTlXzGm8Z2v/2tIuzaGdK3waZza4jiAh
5uN5qOM1h2+Y0pl2DuiZ6vEu4vVJFFZBZdrKtU+/XcsXaUAyqOKFBP+Bs6U8ExwxO+mLLXjhutIc
Zx2Dqc6SjG3/zTa49smoY2DZBbVCn0W7+tfcxqwM+ks164FLqw+uQv90QK3uU35Sh4M3R2wvpJiO
3QIv0CUDn4AmBqkb4yG/NseJ7FzwP1tv/xgs4nrm1Iwhfc596kHP8fCi2bPvsIyUK2+6ThDEXrrN
qqyI+89MLK37BB0MliYqK+/ofrTkp40vj/93RWQj2hG7ztaDgHag4nVXxsqrMSPVT0LICTaTkiiJ
fynFCo6dNqKWS3/RWyT9SgvjNVba0jAPPxEoJQTqEJjc1tgt9cHASQHXMoJRw9tywnUzfNFevZl/
Z/JRxm/H0ze02Qejhx7nqcrCOYxdlEf3WYhz2XV/sSAOOPM3db0qZfmTneSazeK4EVAP0ym7ShNf
BwENwO65Yoj0I1h1elXBw5o/8S8VWUvYALtFRwEhCoZFyeGIBMxpazreAy7e/viib1Goh71oElEw
EfEwervkIJNlmWp1Ft6HCloUfXCYtE4fGJSIIsYKVAXpwIIyMa5KMLJjB1w/hES+VSYqgZWqIjhS
zyfEc50nG/SPY1UrhL1BMqLxhW3NWolwBEF5rAVV1fnujFuOnaQqenwQZSKMJSnIPQJSskIFdeF4
qx5871VbJjpiA/Fa7hn9lDQQ7kHUjoEvqUOktR731fjodEOQZWU+MVfG6ws1OTRRI14GwS0nOvPH
dmW1VXXgBSAXuRK6YGUfnH6SDXPgprdVWmdaobRvjPQaf29M14riEvyPX/KoMO37u+gw+lf7jmss
rAPPuMGD3uTd6qFARmzNm06Ohj3kna4xGlhU1iWMrje6d5P0fav3A30NdHPyh1kM53ejAwIBGUEZ
qWOrdug/oK2TqUvQR7UagST+WEkBLfymrs2hTkEJ7HOAuHqmXZFRE0eLnHCVSLXo9em4nG0x3xAh
NXBBsZsZMbrF9EH3B3f3v/HS9P5atcRIhXRqK76IhGQ05DkyVegz221oKKMxkR4dvd7DWZ3SzY/Y
uDlKE49e26e1iHn5y7c9lo3bxnqK0Zpf7QD+zleum4mFwlDuTxStBUXfW4knAlsRGT9KD1XsUZbx
zU3Epx0yjhpkfj4rUOFzcHROuDbveNg5DDYwzVbc2Gs8vrt7D0f3xGI6YVridtvT88PGMZffvsVl
8WPsamZGY1GrAmVMsyAq1SoC5TnC3yMtX8FxXQnsAxSS5+yX+/+MwxUgYhFn1uS4SxZoBxhCJ/jn
T16Z6s2BpiKD0D7uYuezcPqkwEWtETXvHhOCH2/tl1nx2iBKSCqJMol9Dlppxd4rD8SRU9jI4iiL
xVDZl1rdapo4E0LOGviPYven6cAT8IdsX6v00JrhKJjQaORf24SOuJMd5vgB3elYXEp3UbV5i39C
scNZIuNFchE5IIFXCYtzbH7P43xKgaI/MCjMZRqw24m2/I6fUjLvODzPDpqdTrvhrb2E+jVfgNu0
enor11RBjL5oV4MH1dCzEha59UOZ/nvP+XdAVQr/3Jhbvc941YF552ej+USsP7KV+z00W5xJEAfW
4F7ETsmQKYPaEaHvYRrVzCZuQwaWzIwUvoGMePuaq5ykY9uBQXf8NFiY/vmkqX5/G6cZXkNeAu0R
4V0RPcWsBiyOcRfYtNsyzsP4ZIBxHPa9+8sF4/WARLveBQA5bG7iUhqO7KqLLZ4LLl8WgKB+jVU+
1MtJFMqUDUCgQaDtHCmIfdyHMF5VtnPa+XbLjj0o0cyVvc4Cc1vtuYEJzfBA0pM/Z9Xp4CE58T4G
83BgMsSRNEyneNIjxtgOO/deQgtntumuePphF3u3uJmRIUkHm1HTz4j2OFu7WZ38XUzNmb9zTxmE
P2zuZ+hmX4OXzKgBUejyKCzKsNZn7qggvY3CUwlSInrKZhdeZKeAUpHdQj0EZy0IO1W5WEK27qZ/
RjYCyPj6uNgRnG5mHuc8ygWxRF0DqklRcR4Q/gaUvpKTqRCgzY1UZEQtm2we5lG6XbLSfZMqsFcT
BC4e7VLFvOYBikuyudWZde4KRBWJAxNn/U48RKJuGt0xiKmUfro7bZm22ihYbe9hJ2ikb0PNwSHT
+BVkN+CQc4p7zpsHoyrmpo1udzH/LVAJt1ey49YjTvoZSS43Cce7oImOYW+8PpO4ZYUr73o/Jyl0
EWQgOUKb4VMlahIK944iDOw8ZBGattvpf0nOHc7FAP7BDLMgkdDY+DbZglBJkNO8bP5RlDZf8IZk
4LROJQ0Dry2vVxDV4qfW4KwcNWHza0y9CpSV17m16vVndDmJU8TiETZJJusKQh6uQb02DO4iNYGT
MWp40mdKZTReELz2QEvhEWBc5qM/TsHi0eImh3mXSXDM2/yLAaZd5UQrHYasb9pOy1yeyqMmai4R
MPxJmNS0faEGDSSJqp1GNe84tEzstNJj+6vicHAeGKR95mBvV3nlme03KMZdrbjkhbmtEJ8pT0Vm
AYCWbj3YsSr7vNqE7oxMwGL0uxPiSLNz1Vw07GUYJBL+JQXfGGgiI112oAqnvKFBlc+7xx/yYS1N
LbDbvvKWLWa516EeinUZ9k1XSnAS6ZVbe1vcdW/JTMoqYrV5J3rxypWsk9gtlfT+RTdNP1/dwn7v
eWK9VfZezSKGvOQcN+I+V4+42CHyLDzklCFRT8ZBg0LCf/Wt7WXvA7dg70DunkXgglupU/WaKbR6
P5Rl6gs71W2KniiDdSoIBFU4J1hWcNKCg4Dq+fWVG5VG/lYzZa6yRGldrqD5WfVbWZqkbCjGn0z+
1fc4TuTXLj4j9eREJJHlc5TgcQPx2L3YijTKRvoTp++Hb4t/5dYXDXrs28JzIK0tXkQ7H3yLdnoA
quXmEClLkTJuzuN/aSUb6n4jZb4NywkwqQshLfgKBFNFPr0eA93hzgfuQyuJ6vRXIgRSdmhTicS+
12itsubvpS6QUljfx1BgRRkw+rkyNjjL27Y7XDpw+isQTk10eX8QN106DZWmwZ10OccS7kQHBlPa
LvA2pspXO557AFibrthhxFBxYU8L6dyeH7yLn5cyirUZk8+TpMaEsW5/KS3xegogFQov9tyW/VKL
Q6eQCOFnzik+qhzmk1EOpRjJra+3vKmkAA76TeY0jFKgdOjR+ooZTbiWnK0ZGH1qVIVneNHVBicV
f+3tMkT6xfATNJpsJIK02BUKidVypWPIMDEpTvQ+sE5zh+Sb0hJA/P/KOsL+VZ437kbNLOBFR5CE
mfuRF6bTmiwPipSNBfLNhfQAy+f/0YEg2d+KrVhV/zXYqmNQ5/YY6pGvK2TtTN1RGe2R23xyVFx0
CefL/ht0d+7luRDUjcNjYXYMzVfuOPOHm4SJpQIgP4AHPNZxM1W1Wgt40xpfPvgS9ry1ORMTJz8Y
nvjvAvsCSO08ED3eXlKwze4gqAbngiLBGk7G0RXtK7sk5G/6+7NJBqadFqN0l7vNmajMqszLi1RP
4U3wUHyOK7xHbMtpJiABCsTniayqGR+yXHvjrWa6wXPnnD9wpjn5vvTCUV4507SVx25lA6CbxxWG
dJLun2GlcoC8J3ZDHskliVXs59SEx+vkZ5SRFylgYmFvVsAc7/fvuDticXnB5f1c3XqIg9N82lzp
0S18tzF9R+SUGxohpkvvhK1mkLUFv/a9Gtk2NwO9ioMVdS09WMx4s5JBnsim/S6oXNTDIzNKX6bd
vTBNTs0YEFywLznhPuNtQtlq0PX6Z5lrRdaSOap1+/64P8ifbt7yu9HQLCT1y++njN/Q/yRbwRM0
vMyRpdHpBtAdMxcRfo4ceo1ImfYR1W9JiFMJ1EDEGGzBrzYb67qiudmmwTUDaEBhWPWu2DpurydX
0UKCPgK8mJnggqIaaCwemiIcd7wj8vX+73vVqvZza942iRL2PpvQbpbw1wX0Tct4L76MzxFcQMSo
gbh4sW+cHHoLFFaRCC3mBW8K+eC7lrE8WdC5iSJwin8jyp/NazTEysfCiFalc0n+j2SmL0Qc8czY
a3moOzzWc5U/jdpIty0ZOR50BBYa/yDUOacbjru/JDJsxKM4uJz3AL1p62aw4YwSnBcsqOQlpF/w
MJssRmNaAp4svT6yRorEoJoTS4AH8FmZDEqGiRGApjn7WDxZEh91hhiX957xf2iRm0gsmNcD133y
eXZLcn9yxOU3aiFpJCLAlrFy62YflHilzUZCwmMZCmwxREpYFFFPsEN/UC0DISIDmHYcIOKGbfrE
6AsMVwZ+w0jRd/bi+aj8kdcsbWcM0axq2WTLMxWMI04ZNazVROJL7n7jWfe9yUwk89Rp/ssa8vmz
5SCgylsubs+vqGiT/r4f41SSvBp4YjOh2b7pC5EQIqyg7nb+v60kQP+atv2k4xxrsmGULa49oKod
+Sj+o19Bg25Ir13cyLxevJez+hUQz5BY3pkaV/K++H/++Vnt91Gy/EpY7gKPekgERl2Q1G60kzJ9
HIGXg401wy6ZCi/HPqufucjA6X/oGevPNI9EJkxKm8FgwKOjq/lw6ZZE62ZmnD1PS2p50i7a5DsB
y1ZGpOsLL7Yp0+KgmePZ9o6l+/Bl4JN0J8Afhig6l+sSRoUtR4pbEX2P0BPohyv6Twy0h19M69xB
pglkuKSkDzBaKse9h9FTJMwHRwes65XINzcMxIXyKCAKqVbnN4RVMXh93nzbEIVMHtXXK5xFq6O2
bS2tFKuN9egykabKHDR+eN8/f0zt47hUt0GGe0swUYCm9ucySqmDEe/sXrYPpT2sRbxHxx6klJPb
edBPS2/lki+dS7UGr4cNqgeL6Ruvqi/W8s1w+CzcGpjaSvf+RFESwRMgQuhrGZhsEAwthwryPqDT
9O5JVhidVOOdI0O+zdaS5BSbnjDICIoqBugMxIxcm70efW5fI+LGNDnC4VeMHehRx+papo+iDTO0
RbMK1P5dzn8QIn5w/pvwb/ki/D6yuVCacPKe04dJgBO9+lml3HL8gHtXyak4blxTbdvPyPOi+Sqf
NgXNGv8rJrwUW7/8nfpplp6m1bCu583x8OeSP9I38vB1DxmAsOk/EOc2r/PQXJFbY26aEsHFjnFQ
q9maBVOD0byA4ghi0QQDtoUPFRvgAx6+QpPKM9d0dGZHtUpqZODT8wb4Nu05AsaPQB0ux2m9jlbA
Z8m0BRNgNsaj24/YguX03kRtSP/hqcSG9All/wdYZggY3BdiwrE03VAVnMJp8tcIbV1gfCdukyqK
atezGZ24ppfR7/IotTgIqv9GTyq7JJa3JApekYOTftKXkyULGZvbKf95tHDRKqFi8cVHsO/VafOA
P3qopQPEDg/WNJpIq3wSqQQABvcOkROP4wA/DCCb9p2NAQ4HL3jOUc/8euF3CRmxgIEi7icCqv6E
plAKg746d72mNfKPW0Xdd8a/qmwQ9oobbtfrbCWF2UsFKU0G3ErqvhLecwUDW59n4A7rswAnB605
E/8sucDAtDPrFTyAIeg/lzTBqKs691v6wZhyGYL0v3vl9z4cceHWO4Q6drQQCnY+70LUDIIEIhxY
koflqGtfpZEtXsvA539th3vr5Qf2gAUitI9S+TpHDTN8rZpOMOhmWus7eJL5WY1RT5JA0HwDiygz
c5XdramtFJZs8aKEFauR0SlhE/dLtyxStaSpjmkKDDYdH8t+HOCBAYcGxHU1HOsU9Sjx4hPYP4Nv
OeI2MM6OAoE9/wpdbb2/B1/3tdUk309/uqghZZU+uxdKdTUhPzsC+rmaXSknuS174/5y16thtx/h
bx1d87IKsUVexVjIozfdoyUX0TNLi4RHq7XQudmJED+5WoAX3nExmXb+sFkwJAVXv5ZWheeAIKU/
ejCHJz4rofV0MmdbVkBbO/fHy55s0tI32bhfbu6Aawsx+c65Jc/MwPbRXo2G2EC6YgTwk4D5elRg
Xf2e6RoOn0VpCzKtfWp2n01kZPAhAzuKS6DnDRLlAIJjb26mn2Y2RjevXbSePnyTGDl9XO7WNQ+c
9rlA9MY/e/NLvUMmb3lFR7BSvXwckfhbN7bgwlPeBXm8102d3hmQ0PQPHTRqPDBKWSr17Tm+u2mT
lGzeViTyZJSn/N9MdRoJuSzC9GOoUWYlf1YpcIY7U4smh8auR8pRj5xHHeWPUCUZPmosGz1Pu13G
H/VUpLC+Q9+1q+/jdSVPibSpI9TBiAXxfKNVJEnCJ2ClXAKUvHMsohmZDEowMlqyzjfBdFqkzoae
XfjdELBAtFX95uH45iuD76xRU5nFShxcVxSRrXNC0u9gg4wkj3DM31qyiFgSKLM4auiYXNqpvcJP
jJq5BrO1k4v0yuW9bpr0Y77jCtwQq26myvInT+wD0CwWnw9E3Y8prjdNA8fU7Za2B/kCywk2jHmP
uRrJmFSwzYkGprvgsTVmH2cUkDrB+8int+x00/3NOxemuMwK2rQFvR6U76aAwL+6fL92lauRi6sH
VKz/JhKq+AVWnSRsQfEy8PsObAlVCwFypy5isAFTFqgDODqeJ9mXK5bHNq2eEbqv29765kPilK10
7/qSwjpfM7hGw+8tJb0soY+MBYrfQopxCv0Jmjv6DEhJm2na3NrVb7qaG0LMhtoWWQ2ac3bMUl2A
kdJ/IABn4mQ0gU6DRIj7Zhuld9i+98cmJsgbH4JCmRIr4jjipmfbH+W65BXmysmTNRnP42seH1Dp
sE39rjoPgiDB7hf9/yPjgr+P4RxyR9pl/bW1Kz2f2TFCTAIUsMWNP/dM3PTvUU6DRvEIhyBGOKRQ
UHxcYMQepy7lVi3RR/m6DEgU1HV3t6NCUCPGE9HAhs7tfWFdhGOMrgD3wY20hkzD1Lw07S5+iU4x
2KPbSACCREelqCRD5QgEz+5I0sGDIemEKUVOJ+kHnDH104EXH+fIUBcdrJDKSJ6GVM5c9xltGUhZ
Eo6S1uUwxQkbxUUN8cIG4zjYSQVefdSNVyYiCw3kjtavLq+ulm14OUmJ0Yi/dks9zhWufdmEmZm3
8gxo+jRNAhwC8ciBwBG8k80crEtYIW0bLbxFAdrZqeNNa3TQVrRb2nJ3MsFEeAYxFmM6bWitV3gw
CqW+vP8K8ze0oF9E2KB8JWXhZ9s8P5WjzXQlbuFK/LVCV7j9Hn2lcp0X/1HwbUWar9CMQn6MOaGe
3jgxCPd2r6bHEHPpskxFTKOouoFXjnI3zSmE21KZ5DAYizQpel7//AofL1aK88V8wWkcn+zOTuXJ
N+XLhcAdy7woS4iitjZhLc4XYq4yR39klR/+jGAwq+nuf0hfV3xfmrBoA5Jbv8pmtRDxRGZ2+kCZ
YQXHa1JxIhaVXH07WcbDUzn1lkOZIQvyUt5xmljCHyGyOj8WqWhOD18upE+T10e15gBKD9mFqIGf
EgmhPWdfJeICLHFWhCKBuFjA15jYLQh9/Lsoq2KsOKBc9Xol4WElrkXmrto45G2GRaAThTJQ3iz9
YONhsqa7s601sINkOOKVeqYLPUTZYzM4FM0HegiCSYp1ZHbZhjRclTROaIv5jJ0gmgwhIM3Fgfx9
NLI4P/cAYxTiqTXleMXvUeZLgW0fH4q5hFBODQqXkiTXaELXgbIva/T+90TrpnWO4vTyJTXCu4T/
M9nf/2zF42r+fYd0m9qd5gChXICBESQ6UY+Rf1rXtdQ4ziJcvxXjo6HkVRcjDAf4Cow17ezyTsdB
AxdEOKr8RF+y4HeAh+bA/Wcjfe1VaBrlD/FV4UPK5Z7m+3OIB0wjbdQKqaAjPASZfN9v9ObDyiUc
xAb+QI0ngbZ8CgjA72CdCCXr2/Ux3wtML5FJbPIeriZ6BNv9+7z2LoWR/X8Gs70UdykMirAQ9ujz
jTO/tVnzsBNl/kExH+DCdqg3itXqxXZa/PU/1fGz+tvKGkh/1nttvmNlJWOlxZdT5L4pAs6wVmYj
Nn9IrW7BX7msu/WNrFJ/WFfXFxmAYUGJIMFksWWVS5hOeTwfnWZSCKyd1t381XbMwcb8y4OX+5bS
BwqW62ygvXyR1h6fKRrAnGj63Fc78kEdzSvLM2QJGLbGLWNNVX3AdPqeEg3WsovDSJlfjsEOUaDl
5f/gsGIh1mfDFeWMaRXBqnuDIncpbw5N9+4Ux5339E0OpcXg7VZfOz9u5wSEvcZi5xm1gShB+NAW
W1FVBKXNr1qEofdwS+Mi6V7sIYDDTD+go7z64fZqxXWBRNts+pgZSuhHDOPpf6APjKfqn1iYFp15
kkpgSP83Y/uv2AOMRoJOFLKxMR5vtuzCShWkOCnOi2CrxeCagtTW8W8h0lrVKm7F1AWumlAIVOgD
k18NY80XCyR5+8M7Va3UdgXTjxjAgYTwcG2VFtgMpHgZbLc8okzQlXTMufi3Ov4BpbO2lRn7VAzE
ASswwNbwOE30u50XIfpls6qeRdO21G/V37N7jyiGCwzGDDwiGBa06TvAkMJylXaM6FJdW4Vk7Lwb
RraYdTJ8654GwOf5W+Upd+vvvizfmWQtJ6g8huyaRGARXsavBDoHoq6ti71JIC4EhwjSd8Y9qlBE
8yeVPuoPuxzx2QGDZ0RF79LGXBwdo17LAnIqnTFEnuxGUhGWE28ZWZnbQ3KfVqqPgbwCZWC+uEDZ
84CVe9je9X6SlxTGL3WYsF+rPf198b29RXQGKhUSrW1CKCYiWm4xfu0WIdGY++kSCJb7LpaFEBqF
gVY/5DW2zfIhPzGqCMnAZQvgUeLRoBF779iU2m5M0P4frpbk53lScQI6BT3xLGIsV/f/Dcy0XzDS
7Ma8hkhX88IY0Bcnhgg+g28hi0E9KlqaH4KJdvt+eKx2dkatzrLIpve06WuaMYH6ZZ7xjuy4+fNa
6WGR0E3mBLiPaQnIKzDKTjt7K/fvmbuUSAQ5iTeKqnL4xRdq884FzcKoFOqS0fIrDaofMW38RUZq
LdAs+l+1Kq2N3TOO1BlgAaS4+IT5cIDawXZ0LfiNTIhCo71Zps2i5R/asW1jkV7XZeES1h/3UeeN
D1Uk2rZYAarKMounOb9kEtgYtZvqPgtCTmjGlb7JCpHJWwD3mBhSpvsIBXOJN/DThdpmYV8GzjIq
bxwmQBSOBdjVmG+FFEXBOiEZXAVVSqnLkTDP/endxIx9CWn8h4Pu4LQ3P1HuIpWmHc5cIFDQkimn
nUK7ygH2l+U9mQKNS/YUCxzY9nTmXc0n0jc+gJO3rsOo+H1ZeHA9DPtsVEnPFZXqnrdlErUgiHPV
y2Vbn3ot9EIcUyRdgz8fYm002Wczf9FG345VMRJ+SqccqwHKp0MVyHzXdmGThrdmpxCMnprurJ5B
zl8ifr+Yk4yG+j+QUX9UF4Ym3Bvlkyz1XyuKFoNtMObt7Iccgbef+Xy8fB31DrFJe9seFsE3to3b
CkjEUWv79sYnzJ6g3QLwoEqXlrW2FMj90127Wez4o+dvt4IZDvpDgywot601yaFEFeT3P1JwJucX
rId0J0wSuBembDto9UMqYRxF9R0xeyM1AT21440UH87hQvrCKDZNT3hD+NmrV8fBQOTGLl/fkqr8
dh2DO+Pp/gqsdvmmZ8OHqhJWmX3iLvSBVF03RZKs6ayMTuaCCUvmnyOKT2iUKVLBjotAbRdJimO5
N9NaIWiedOn5USUdpixD7apd2K3JOL4pAn2d6fVxeaJCQv6D0eF9C46ubYFJgffYleshho+fnYor
w1JIOSe1r4lhPNkSruOVI4B9LsmRoxhwDXASea+3AxB/ZKQH3837pPBnE1/D4elyw4dhFQZgIeDL
LejEV8ekeViRM4/jtQEJPobM/REV4BpLvnybNcSjJN9B5Y8J7vA8rOPGuoBhR6nKYSfO5DXe4oXv
h9slfi/QOQG/twF9PEQWYdPvii43FjGm9U/9EcK5kngRgD5/7ncd8qHqHQWWHYC+hbumGqQs5Y2l
v0oiDv8GpVyxlR5GTB63Von9R9f68nnNccl68xR6dIWN99ZXMvTsNzXSM7CoXeiJ4O3ASdth60kd
3n4qHvZAwrFH+VOL8Hou833Fbazr/H1uqbhDQPyAhZHQcBmIoUkqGFHb5GQkaXZYSjn2xmgGGX4q
CYPOGKZWS/o8asAlh83tg1vceHo3Vwxy3ZmPKieK9zMP72JVACVnEQ9ZfrnAoS1sB8+Y4J7nSwOQ
TG73yUEZZwqADmZzNh6jvDIm+UFpsOh3cbR3pRvM0gVuzd2hz5W0+6ggdZ7AmzNVNFP3maDFPJlc
akH2qYZsxi0jGUOvvGAY/kd/WC6fVn3/7Kwh8eu4o0k+GusKpQSREZZNja+Q/FGG7aoI6f77lkT2
RGGIms7e4E2Nsqd1AlMBGYDvjuUPJapu9cdnRpAv7jC+ksdLJJ8xjKXGtZL43bFRPNSWqUQiCmhF
4QBoF0zzjroDWMSeDq+cKI7jTYYcQ/mQjwluAZVAJSqg3ZZforfYoMBKszTeEiV5p1dG340X6/Dt
bVFo3wHxvrg1rDVHCa1W4xwjGD1Osb30X++h36Ai4WWOT8soofmM1ABzPo4kKiTllq1xuz7nRnon
2TwHM5htJK5lQ1eiyTkpOSyGMaZEsTUGq0cJXrYbbY9ZmUG26cCIm5HjiO0NiIqPIOb1KUr7MiCE
qFAO/3pE/HfeAlqaUP4HU1TriEReiWMZqzm2vM3zQVG5J5OiiAKUR+1njVvFlZZIRADjAZxYnwnw
VVUyeIKe5W0fxLcAhq0EqLBfjd+F/dMa7e7yk+zLKeyC2GPes53qc0VUA0f5vz5BhZP/QoFTGbgf
qfaOr4l54WlxUtNRmmVxCu9GTik7nc1p4dnqwh7pGJmyNoTu06GS4QokS3sJKQ2oT1+OTr1FHtP4
NBY2o9rZiLli8l5c0Moi0qroQ+wnehlTRYi4+m1pAeqxRHYIlgHicQxglYNQAGP3HhbviKm1g74W
Oh81Ap2eqt0yaHaGtoAypo925qicMiYhpeSCywFUk0Q2X+wczNQedLXZ+1q/XEyTb+EXt9Znz4Yc
PA3yOvPh9iXLgdZim8zKymatDPit5K0rtcSupM7yf6f2rbfh1AVNya0rW/A6JEBElhFzqnPHTB6V
QfTq6tOqQiGlrRxVXbFWZ6ZbUyUVxLCAFRRNxW6eIaxdl2GZ9/Y7Ry5q5T13doykL24/cuFDmx0S
E5XBxzE+DhAfdeXVrHJftTJIjZPnhuvZnjXwt0uIcAxhDokbH5FHPFXS3vm3i0NmTo0MPUq5wOEe
Cf2d8ErdE5wCXPcfg3Z2r8hPeYGKBzWYJcpgVRzdpYto2D+msJnzvUh7u4CqR+8jxSdyEXy0JdYi
g0ouznei5/I6fNMVq6rE3pF25z0Ol51reBeNIqdUlK724qx9XjO68QgwoBbTeYdZGOV7FtFSmdky
yAXi5B3CuKlwmKDnxUywP+kaCBZNq8oRtUPlvLjkV8C3vXKjTwCPZTLgJj2eOlR1UjzknXuFVkwy
kwoKivGKr7qXQgSvp11wLjHF8P0+N+UhdQCsly17l48SUoMYLkVBD6G88MkLSIA6cb7UPBtRoVjX
oWZBcmw4gUBhlyoG6T5GsyBVoBVWPXSvsdH+xlqxtUuM1cNJNcgtZw5tHFYqM4ELDy6cGtC+cvR6
CXcEwohatO8tQCDpeStDnw858mHxspBams0CLgyA5PlU03uKqRaEccdLXzpn6NTzCZLZjlZhIfG0
HPX2/eaOzplv6dLDgsoHe+/oiiWBNddcop8Zza9DJaWhQWooTmSuaqglh07bW8PBlOpXM3ILt1vC
IYBLdj4uXqcmQ/jqpFa9F8VvhImDcLMSHn4DY7CXhaCI0kyt8qphavKjHiqoCoQHr4sGtXVxh4gR
7vEHAAUrpWS64Nqw2gFMVZnz+R+H0OdZJi7teYvJo3H20AxzWILJKdfB107muOegFM7ooam0Sfya
eAg6iK+Tfn1EJvfyxprIsWu9xOHXJCDwsYo/3kqQLMkMpfEAaHpWRfcScdwt79wKTPkXK3b4w6JL
5JWYIFzw1shom2SPVEy2mLEijdf852R/3YUuRS6SVyq5UW/DmPQk2oBo8LqeLopCber0QHppnW5O
owHzU9FLZZjhJkYVnS/K9yNuL5lzT9HeMpVb6mCMpZAht/vzlXvY/+XkHPF6A7QHOo7KuzVvkEer
QpaFOXJm3Me6Nkr26dMheutsSNg4uEPmVSFTj37HMVVbIv6khNf/kBeISN5msYJbh/0Wwl2VZ91o
KJMdTW33Euoeqci5r2k+gqBbsvJjMjv2dxcZI9TB2dU/9f7j53PvoGT/mtgachX8/Z+vbYdapr7b
iVJJYMfSrhD0/2E6Ml05qW8lNBYRsyCuMUcEsEk6M6LSu3G5Yxnvok78MvKZ9HyeNlZD3BwzSv0x
aBpoDXtIIcL2tnp81Utw18OENVUbIhbTWEoRegPC/gu2TFMgjx6vz858qQ3cb2IYxB+3ZcRDlt6a
jQkWuJHUo7+T65T2aThZV96NsqZscJg3vtzqSVYw/Adt5QVepks4/4jsz7ol3IZlivgffxzX5qNT
OJ1XmztdBNj8eh7a85mJpLDuVP+gYc7LH+MB+mXO3A3tU+Vm4lD8mcrdu2UZXfmBarRhjUXe+WcZ
SY39EmsEegLPyKoRQnnM/aOjfhjtzaMNaZ4HKXr3bYUFhutoS8uk+8XIGPTSiEdcm15ijK1YvdnN
4uev9cTmq6/d8zQKLU/nK1lP3z3SUTmZrB1qUTyepwSPvj3kcxy3UQLyUMEEwN8yjHRHKs378y6s
NS8pn52lXW9ht7qHU4LxyG4Ym/YCBMKD2aigHPbhivwg8Ts5BCT4RjlfLtM2JgxzFi24FovIlGIW
tnXeYCWm0sn+zbJtS8q5/mnSKeuvWUz+U4E1xPKL81PTL5fpapgN+oHZix8u5L1BkMvLV7gudKcl
xtKIrsFMluv3b2RA6Kmat1Bjg7tLWCXyyt9Hr8RgfK8pCO2LIhysStRTckU7eUcZpcV9/ghPh3oc
MJntuB7ot+3tIiZ212Xmo7k+sz2z/QPxznvmO+frV/qKF3UnXSi6edANnenQc+v3ELDYUJVUDG6g
39cddEAsuFUUq1R9J98fHOmMbztyYEz3ikrCYiv87qPwg0asfGpya1BfV8hESk+ON5hUlzfXPgDF
LqAxHohXgoi3n09euGErkDHzzhB9lCtSHrkmVN4pTjBKy0ZpprjL1yHhsQEWoJ/AZuB7kWfDTDc4
VBGKdQ4USBs5VA1Z9PpHc5x7zdzG5YC9iThhcCbLh+2rMhAX8zY0sN4wmpl/WDeDXprEN9PzAYYw
QkuA77DKe4UzKxjuwHBNtV/Xp1Qhws9NqEZtf+JNDW6wEx1IGLDVP7UdXH1DPFmiT7SaRFHO+Q6i
vLmG4o7gLj7RkMUxb/VZ3HQmHlHoNvTjFZhTuyhO6EmhlVVttOYBRrdBlQjDx9axGEvPCONhGjNh
c3rHxoi2ZX2ew9oKuM9BX+L34ckmjcKc+YtpGQaMpJ+2YSTbqQ09JnWnqFDcctFHLCCr2yEU1t72
akz0xBpR5bWcRUvRV6qidcOnLhm+a6mCGI+lm3MH16mSqZOc6sPX1vemxcA+nWVKLqpyYHM8bLi2
In3BSAa/x823A9jiojPS4aL7H+sZjLmWtVg/FKcp86R9o4gA2j+W7D24LPvGgLxSG4y6dWjnQPN8
+B7ym0Gwxs1//xdLr9bv0q5zneh38LUxs+l1vhbaARzWNmKD4H84D/XUThjZJE72GJbGlZHQIVHh
JShYWU0HQDOcrlnJR6B5twEB6TRAkK2l2trUN6WjAFIU8foTPz8/+X5VLsRrrWlWboz93ABNjio+
RZND9waBhQRIJVX7kodqLeDPbSb294vhZauknr0S25yM+/Rz2y62hRKFfRltzZ73zYxEcY+by5mz
73sIgZwVrnrWBdh9h+D6rpIp5fLGg8/bwH0h1hUHvz4DTb1D6ZeKM6uUWLv3RA6naDAYQvD59yla
zWHmi+OBqqbuMJEyi6p6vjHhaWhPlUwtQG1BgRHLu1sThJXUOsJEzXXT5sfWpnqwZInHLSXKwGxy
1nA0KaObITqq3VmVM9WRTWn/8DSu645KoBZAwL25HdFKvksxVScmjgpRWoloK4Fs3oSVYB7/OcmZ
ZxrvoVYf1IY8JJ7Eosu8Hfm9OzHgKk+wDvXsTyXyXAyHt9R8+TWp1g1QBqIouq2dr9Hrt3tuA66D
EBBYPdrZO0RvvBakozWDwxGNIz0SfQgRVzifF4N0Ccwf3KjvR2SEM2PqYIIfntnBVM4SKgx9xNGN
+XrxRi6TFbyzhqMGE7vLZtiJpUUuGCHm6AjPU71FgrhdGEWcUzBE/lGAenfIG47JwplKEJyZ8KDA
JCe1NHTcE3BotTvFsrxHyKspmfMezVWAoAx32/dxKpNEH4c2RP8Yr3eL6I6XPJJ1F4KQnB8p1FUL
nJhVzD9YB0y4GSwmD4Y4z6lMOsNDBXERhMbs5Ei9ioEEkHKT2aBb7er4jqyZCcS4EAtiJ/agAE58
cf2Xki6hhS7MYaLSTaZYZJ/T5KjP18ipKqJGY1CR+VR17v7RWHURfYJmN59qunEgUfpndgnVvB7q
V6Nke7K641g+khB1zBeT1/1x9oIK4pX5TNPg2i4l1M4z+OaUj3CGoKvbWdBbQPIrPymW9wrWlgJE
cwLC117zA+A3M4c9fEpmQ0GM8nkcFL1cFeSh2lMh9H3UXjkjjmc62ejm893960lTk9E7Hp6Vl9f7
tLZf+K496z8vkhIo07CL8ZVVteFtcYwAS1iNpA2EJXInBxYYoLgwQlKzibpqgtxB4jJ2GRWXmaJh
hZ5j+QLrfC7F5BSRPjwl0pm5E5gVGUU6ADdPYFih75lkFxJPgO2qfSsenzWmU4PDRHeEPXSZkPKb
ngTT6yEEHbVEqnjjDHLrZ4It03vtvPxVfjUDVXEDBInuN5woDYU9KAzTlHr4H8x5TuJv/taKha70
sfcclLGSlkxpXzUFHyi2J5SB9Zc2GpqwUkQ4k8107OwIE8VOMlPvGDt9Vru/r54vbMbPfCrNYCLN
4kSsiOSKD/H23hZw12cfL6BqqSo3ZYZ9Z4D74CL/T8raVRGqLYoRpd3VW7kqkyfHxNIkaiBncXj3
zWYttla4acvAT53q6CZohlP75GUmWmgPxBkVo9agTjHDZ4pQdmofNFLh0r8rOz0ZJc+i34H0xVbM
AFWIhEiMO3Tp8vBq8WdFXWuVmRwwa0h9BkZM28OG5LPpNqlSPGK+4F73JqTXfRvAoT2esn5xa6/K
309+CejtXsBeOmylgIbQJn2LyikcTMs+QT/x45m4i9KFwtuZxivhQMISmEwl1LQTC1QdyeuhI+RE
2QZ8vIYntNZOzsZk0t6KriP8O8BFyUENvvyiavX/U5ZijkMal3HIvIssvQmND9wW/vp9LwjQO8Kr
ukFDacM2x/itmN8g9HiR7lemYY/BLA9AH/4VGS/wy3n+y3yYwVujQyob4m0wJN8W9DEHChzIkPMU
d08XVh8L8fduuCgtnaPODwXxINd/1tDem9W9/gobXNDwK/FRrcO0FGj0py98qHA5WY0C2Y2wfI3Z
h7H1zYZh/+gy4M46Cp4YauxOg8t2UsT9SMyoaSHXZTrFivIqIoJJDcn9ClAKOyU6BcuADfNlrWx8
VmRX5NXCWDtMMLfOn4+5foKrCF713gJwoyvTdQMSMTDu0bHNmfltV/ALfAH0R2mfX5bO9CZoW735
zoVHYAlNmsDaUWrGMwsq9Czd2Q8Z6SpWGTMbDYJrbzL7QFahiIp7EYHxoZTkvps2rdzqwUDNyR8N
lpnz8PIxyB479VrWGCes3rUT+tK9Zszs29BZKawWHiNWkGnyITkzDQE8EJltSbZXW8tBOvnpr8oc
bHMKdSlmFhUpT6Q39o7NRQM5CZc8rcnuoltMJmDS2b1iAdiplEOs3lMZMLo8cTh66p4m3MucuOQg
acFBq5S3Qpf8jo9b/BLExIO1WYlqWYJAwyscaJ10xrRwt7JQSlnmmlTn8Z4Gj5Yce+9azeaKEQcG
KSfooyi7axMhUBTL6fQ/2VXdgpE1lXLA4J46xWsCv9q1J6wPwVi89Eqn4tO9WxR+p4EwqHia4qB3
HABm4Y5TX4oPB91+qlFVLf5KbMLeaMQj3BQ7cpr45rAVfI8DmuLhNXUPd1zUcS2UJ6M6AfKh/pp5
e2vIv9HNLrx+J6n5zSSkq+Q9W/JY66dEXlD2EMzFHMENokmvlU3MnWqZNI8aGicdx/3nlRZ4qJ+j
aDfpQdm1KcFy//ChEw9bw4b2tfESoxLeiEF//o5tGvOngXRBZNbXRQXJE+rkdPx+wV1O7TT5ho4f
AOVKoUSBPwkvaFjJ/l3nPrLCpnYGamZIG0dFrsFbwToDeFNQYU0eFwkhanCu41zkflrudocpZhLW
4HBEHcURtnENgMOdLGZFwM1vIDNiga3+hhDlDaYPrr0k+FXDZByfrDbK5sWpwGV12v0ZH0NI5W7j
ToSaYNtMqpXaLTCPckAPB55g1Wk2UBTZ0Ddq485PKkuuYOMM2JJDtWqCxrEbaakGVgdkQRSFOmI2
qWirU6axZf/gv4v/2Dzz3q/OpM+ZBZMTYJCRG2f2l+OpNrTaLnYX0w+2UAeanKMyTnCWx6ocoeCC
XO5hb2SbcuJtM45HEFzATVv5QHQHofuwcdxIJ9M3/3strHcpOEu5y6R3F8sjtC0g3M99zEltTACV
XEtqM+Pk8+ssgDQ9lgetUQ9ShigXAtlY6i9AaXFJRPlmo9at7zgE3YYmbHOTpCU9HRKO9FJ0BxCc
OnNM6sE80T5uMoSmIYqEQ9rE0xvph3pSxTV6khcCICs78f3rNKFNyKWgpN/ldbj+f0jyNB/Gloyn
on42Uy+OavJhUiQGWE6d+WpEv47/qU0s705M80VlfZG5MBpYfJL/tAIOtvooHkvuQpyfmGzO/uvk
JISoJcooV4TAbRY/ta3QPHk/0EPfZljjIg7gTpdqLth2/7ydagVAY+wrshIRQb5Y7Umz0ycMY8kY
jT60gfN58gZ+V2qvrZqWdh/7a1Mq6B6bg1Ik4F7stly2PRB8naUQgHaqiKjAeSr0zMJ0WqoISbej
pUYSsesWMEgCJRFcnCnZojVggufViyJZI2cDmLlUtLy0FzPxjaDejfszvzPu1qQehAd9TdksoqN/
XUIxnGMYwTdz22jkW8WnK7Sr5p1KOZTpftLg0Ly0TNB2w0ddat1GL6Xwoo0kyc9ON0XDNH+xmu+v
a8vcdYIg7U2TmKavhc+suWoivfK7kHb0danEDoEaBK1nqIbkDWVEP9JACQOXnE3YEdrRBMtBet7+
EqVbnGiz/DPHfq5+fZ7RKZ6xHKy+6H2KsT91bD9uzQylS8pr7l12DuESJgHdC8y7aAkWBt7b28z7
lmQC2ES8ec1+XOCFRDIC5fAJblxI4F2J0/TM5LEy9ujFqTFB2OJwE9DL9e5HK6JHDRJwSL5Xbj//
4FUxOCGkVIqp8PMvN9XUdRz7xnFTv3aKzIbmfDSGEnk3gsKIr9t/ZxpSGbkEzMLji/PHZh9sy6h5
Z3RoW6Nb5wpoXxIXsy+KaU1KGfTTtInkJvnRugGoFUfxQ7uoMFMHKrywadJkXPE9XRtK4q2oG6MD
HqltbHXQ/HSu/ZfZFT3sU1u02kSRXAzQkPkwpV+OvhcKJKHkzG5c5/XNN6nIJLumv/kbFHIxzn9I
qR7CgcPMz7MdZyvCF+Taca1/5KJiSsiBPmOoXDT3eKrqy3/CazITAhQpVTeAJjFDSuY77A0YgnXC
WTbuAaP59vlFfeJYdPpjXXS08bqVSVbYZmWQhPRyscaQvjQHSroucCWA4AmxSYBtdjqlu4+/97xu
HflU2ma7M3KYNPFOVGlwPA1EhCf8cNt7P82b9q4cRn4rDFZR2W7C7//8GGgdxFvalEV7CCq5vp3g
zRhcr537H/Gp39pmEGV0Gm/8a3SoJS4413vADdr6+UpvtVPD527mgKzC+Af0nzXy1h04boDScBmr
Lr6LjGwW+CJdzh3aeC7mh6EBZjnxXgoVXxgHq0zz7y7IYWapnIdq5AkjkdsnEmtpGv62P0QGzxZa
G/pP1ZUBsiUQ1rxDlxqvfM+88opZiy7MUi5jELB5EDmrJYGjGRUcNDWyW2uYZlPXHp9+hWLShSjD
ACVR/Azn6NWG/a0M3rX6f6jPkjSG5enxD35k0iKafe17Y3oG5r4Qsn2KBVGAaH0bVDsLnOvHx5E3
yHsQxviKrnqteoV1yZaXPbVBQkAdfZ+x1PwaMt8Sd9+bAccOCo9J4DW9XX1iXiBqJuyuR8ai2P5l
DO2Vk+PV1FQ2PuGPXOX7tteEboPUEQZljMo+6oz1wYZryh7NRBJQ2AoWr8Vx5mbZfGdpTkQaZMYg
fQZNymfKQSJryQP0kcMMDrX9oDwhYzanKmD2thU9XbwByskMuO4auFXE3PvVnpwivCbyxEQVUTHR
lA3hUyt5whiDUgw+7dwFXWaiNm+84AmO0LZuQhj9a9tMA7GgAbx89i8/NeJsPxW2RHRi0p9eM31A
TyqEBfKGdDIBbyZvC4US2S3cYiLjOJ7T+OMzoNm9+2m4AfZy4CdzMVj61Mdl0N3IMVTsuhqu3IrN
ZLQ+3/okQXtCK6uvtSf8ZJvdnuOFINKdpCIn00B43s1+Njm0+EJ3DgOXWotaYfvBgaIGTmh1ZpR+
fKdlJiwttAwsMCMK/rcxk1MfbV/WOjLnbjwKDVPV1pQdV/FLWKmqf/N7lzELfhHDZQBMkNxYkKNn
QIf955pkYLVhAWMHv/IZ0gJY/eJYCADsBo8I7ONIemtFa+Af4jA1yccJzZ9sQ792hgxzP9N+1mLi
GjkmdjkIza6pcIs8DktgeGHN4h5sIgQf7xYdC4gNjoHNzMznQgczZgeBoPWc/O/wYLyqQYtrWT87
kW4/4FHsWhRWkDyGSNp3pFYerdILmKlgwoqeUfowaHQWQpEltxZYS412N7XT7MqYQNZastlGa342
IjKh0cXODRvdJN9Y9s6RaG0mi/dB6HPgQ84TJKHOwDzPOmA8cqQ94fc5ctWP/RiPfYO77MllUF7+
unzdsxSUOvO1N6/jdleaUPSrmJc8iGDkY+RGhK7Am0W2AMZHiwi3SiWA525CaKi7T6EwgXFfWKR7
Hml8nLjFEpnpHfxHxzZ5/XZyCm6JoHzuZxNYdv33C3TgPJrK39c1/myLvegIt5F5gYsiYaflUEFN
U8LqTnHsk9LnPQnYzIMf8uBOMYiXKotlI2jIYkgmpssYJTQ/amEmxkVEsts1j7h4hsFujr7JUWQs
t333THA2dgGq2SyBMoPpyEgCyYNG5j5CSrcwuMJLfNqopRW8SBx6q5fhWt/MSS2z9+8Dnmeu+bfc
yAlY7tPVfZKWsBbgh1TqIdAyyqNVzZVwuXAp0qFngj7p7WuezZBln0XSSAh0QDxzEti0bgHJYCxN
HY8ffIamYq7r5Cd6MlyKantHr8IoZF0W/54pd0csZ2d5vuiX+Xd4yGekkA6/hm7yDuC43vjArN1W
Yf9AtzPBR8OKZrNhVtBPGb666hhVsmz9Wqwn18wgC0BmlP2cHucswA6Q0gGZtnc+a/d4EKjxpOOh
O20m62eKT/oijhP3S/vKkxHLgJd211xwciy5WKO9UkXp5ICV9w1bfJP8Is9yd+wARL6DzM6BZvoK
YgUjPfu6MDd7+hB0gfb9F22YYY+DZovlskKLep/vJfpOwXXgAJ7lVdc3+PbfnH+diLHNSyAP68AB
N3gpeyYA0fkMDPFnvTMEr5zjXw37IWDQgfZm9jaVgeb7h0BI9g91gtTFSPFdN+QWDp8XG8/X3tU6
j5xsNkU9VIPV6i3deW6XUlmQf7ON6zHWEgQo34t0U5og+I8fo3oKTKRTxSADeXHL9Mm3hpZjwVt0
fzso7xo6HewGB18WT4fFIaqbNy7lGgkortVH9DI4XJm/UZBID4xnVdOgKnvEvKruRe6bkY4X8ODa
GO23M5zumEDEdTpfG4ry1yA9gt8clodgQYxgqU5HzsmK9lHFyNOsZxn8HR8NIXLfF4HMhPGw44P2
1cPMyXpWne1FdKmAFc/pbve8hgzFAALcoK46V8PZ1ZzqC9s71iSj+czTfPMrcHsPZhJxbLvJdF7+
kqvn4blqqsBwH4bA+BXkTB29LQdPg1KXEfRsND7MpaTHXICAhF39/LZ9f9Wknab1jDY4c+eCOyao
jj+Km2/zI324EzpXnLKiJw5WFITirfcCXMmTs8alzP/N0R267UtKH1XBQ2fZuFQOnTCAjEfpkMe9
fT6T9xaNQivhqo57ZN/K9tminnGkgdKyAbkUpJvb3BSVTwesB/sMMyqAS5SG2q1zMwbZHKJ3Yw5d
DCAG0NWbH3eX+PtE96eV2c3HW6i/J+uUwJRADfjm0ztfUKW8CrzZjb/uUdY40pPF3QkOdEEgk54U
rw34PH8HX5cGPTcPY9YWeAW3D18L4cVO6Ng9KrhW+XONssA2wUWxf1xhB9ssscjKrPQfeCQP0c00
UCPq9OaBuSJH2Ehb6LhJZgOZg6T84U8V5qDnSDwVTYtnXo5OviXMSKteVgfq97rGIVzmX2avIuai
MaLjIypH4bFkQYOnUz3ygJQP6tXrIlwZbNz8zZzEPBbm74Dj/uE6QV6WggLyCX2ovkMjWRxBW2PG
q2mhDu0E0i/VSa6+AhfqzCGT75wpW5QIn94cjuNKk/1eDCB+jrUNaFD1kZ06T04VKKHMRKNhcm6V
i2MWH6YKwBIhqz3mD+ar2oAysqARKcGBy9m7CFZCmMTP0jr2cnEab7zeZj6N46mcKY8ADELw5CcC
9M6up9NTYb54udaHtmk8xPbIzQ5bm+KHlV0hk7RG+U5ElxYXEBbRFX3OswYUR+TM6ZYFEehI0g46
+V/Qp3kKJLvNSbBaannX1imFga4m5LR5tP6xVrTwAzLs+IBwyMo+T8Ggb2ik6+90I/KVgSgyqcIR
fEOMyKKCCAdY4wJx5b06OS7P+cTnSxSava9+FqvEEzzf3BVLlXzeHrWFOOP83x9CLkJfBKfHI6QK
F6GP2XnYwZqBsWzuaH7UTy/Lmmht1kjjHlaqFgCyGF/kzG2L9WW6gHvuV4ak8reVIF5TSr1Xz2+q
q2I19wGSQcBhNY5hvioTJICkljrGr2/FKJj1dfwI9wZXWsrdsj4OtbUeMfGewbN1t/KTh3FcXQKu
h3qe8xwvL89M3gMi++tZmEsCkTiBvUXqee/xo9xgv94fNYNKHUQoYBD9xuSXd/JA5WAzQ/ZpH1cE
blljffAObOc5ZdCzPG6Bd3NTOnRQwDahYl2b/exwtLzOhrMkKwDswSPgx32Hq0bQlnZDT9JpNMkw
WrnjbGbrf4ItrQueGLDBUIpXkJMTEjQmylDprieCRExMs4qi87s5qEwzQEC2qwbSDu+JV+zdkJhD
LE79ukx4KJ4BWQbBKJ7OK6kaPHZapx3KkuVb1D6b0noLiiHn5FxTvar+1p5JTnGRPgRnt/qphVmh
F15waHbkMHGclAfR+80PdG/DbYjvYHCQ6TdQddZCjcPLNs6Kn05j+HxJy+dWBX4ZUu0202kUXccn
UvQGmg5FpE7b70uJwpRHbJeCU/fQ5c4cgEqfAK80+IwV/aDAPswUtee1kABV0pQ97GFUPmKF5R7i
DEUqPp6bnei1AmUJ7Oe/oP4AXdGL/uDkATRyUZ+OTDwk5rNtGK6m4sJpil09GrdtXNqwOncl03OP
A6MO94VYgngNBa6ko1xSAEjtWFvMrk6ZmJlJ+yvK1BZZ87SQOD+v0c60kKt2gvSUnV0gAVK0VWr0
j6KEeMSp+eh2PLFatBdqdpuOzMhSi5tTTv8uZw1UK3GNHupdOcCLajSqD1HAQjfLT6tebU3pUVid
SQYQZboZ4KvGnr4cKyz//kwyDp042ohOaapbO9UOd62+27QOq6WsO0iG2oYj/NSA0FTCt6BPpUd5
HekF2wH15mQmX8yVREjzBcy0YoL6U4W5eSYKaJMAMYxDSmAf2mIMEsOKG/gu35A7ebZiQsqk+Oxt
G0rBFT+YFxpcL5RptschWEbjo4Mjbo3ttPZ4mZer4lLOBhvHl/OV44acfXjEweODILe3uQ9KPi3X
/iBcTUywLzYWgb9nhMV4MU3fnmFRku08lGz9bKLQvr4zFZe3JhMSenzNwE1JKZwtP7ciW7pY+ae+
0LA/uNEUJ/E4ISlQmAGojerGenJbjy0gLQHEBsv5fkFcu2/IWFnkUJsEo1PuE1l+RHdyJBRmGI7c
Onk+8V75APi2M6uhMx9vhUIYhtbQa4Y8Q19IAppJ16kg2g/1o6/DnySsdO5laq0W4eZBfpFoSOQf
xcAa2HyEPh562t3fRE/lDNu2FWYKpaUidxPW9wBmkRlyCQYmj0N1U39n0HsnCo0ryVtl/HCJ4++k
xDmcn1zyMijqQ6UNQ79BHFDbEZ4O3+TATc3xMwYn27yWNxC79LArTQ1+8Kd1vK83WaB4UleLRqrp
A1ycbn7Nz1vaIYB+/ONioOnimejM2p9kf1GnvyEBw4dEIAmVs5KpjYeq4cFZoS+fQtxhDaSxmOyj
pMZA38/qNOITtmeHdJQYolKukdoM3UDP8OQEp1xgZf91svwYScdDPNZymDsErwzq/EZEutY4qIjx
fMpAbXso/imrTt+u/3mCA5vqYBYiDrKfLMwRtcWST4ZNC1Ki8C8ebSDtGEdG91ltSXDRUeo33m26
Q09W+Dasue87/iW6In4FckIOwqUZaGUPm4imKJJKFv6oBejRyKNlUc3nXdHo479FbUOOyDyD8Up5
DAmnrE9lEr3Ou3LApN4+sNucSF3IFRFpyO38ooiNIXWT/wo8NlaWmCr+axiyMekavFpVELS0zxdH
/L0vVyiGfUrBjpnDzD/V/uOLalN0Miq3YbjU//lAtXuJEOJvL7oZ9wh+IoooQ9o7dW8Gab90iS2O
M9UH4hGym/9tvZ5lmGVe8fFesNTb4/A050d4uxUhuWab5Zz5+C8XKCS8M/Fl2v80moWdDRlmTtUT
NNdsOVnWkIhy6IG1jrmhBHDQIEpbQ4lQ6gc5DgICnSiidY+Y2SUehMmrbf79llSdssHWh+VXgoff
obyO2fiO59jzT8BRMiLSRo+DwA2Y+3v9sLT41tI9dBg2gnJ4dnDsciqBRgwZx7t/RMJPsAPIVzb3
Sy3K+XEmrqmYIMLJ0nMl6xReHqFUvtSYvv4XLnCDPtukdYKhkN2p9tWeweTTgAIduB284a4RV4PW
EfGDeDG7kY6gymnWPAnMvBP3ggiOFVQ7rCljscbB11RsaNHSgHGLLFTfZ+GjUUs7CI/6dEhaR9pe
ep//lNgHyzmvUnAXue9Ze9Xnb8DcS5BEcmWSmrORRIkMPOJpmjC7nvCT9R0q25UnJ4NTSFfNJpq3
WhzG3ZzPyR3Fi7F0GQjtZI+Cn+w8xNcngLyGai74Nc0DAVTGE7fYxB3+E/GLQQQQRmBSAUroU9Rz
bhwqlTXefFGfvMThXK907KCCwBYM3qPPWiJLuxdIhTq1FG6sdSE3Jjsr3kPVw8DCX+3TJdhoUfnS
p/dIZFdYzw2D72r5qIVCZisS/qKp2srgSUakpExjcN/VxDmoTmx0YxTCBJUCpoyWsJsyoKuVLj0d
dt1iV6DtYpNTyAXdlX1G5/S/UBW2q8kZV/OpneDFhiVngt7ACUqdTM3zsqQW6lHV1vmQzd5/hZ3b
2lY8wKx28Yzy7UIHIATmsPvFbp6aevkpeIgYAWjZt4+P6XV/cZCru703vIR4In6CEWsUfwHAqvVk
gdMf67hJR4LQaxYvqvMXDayTwJLy4GU0zfe9Hankxt2/PE4J+BnXJcLxKejKYGxtwYROMoYYEq0F
XRZtchiWMuAPjC1kTLojGgh+pi2VY/V2zPgQ/bgzJ8xSgo4oJP3NIK+WCPxTaC/NRlTzli7rIIj8
glsLFRDm31m0pewiqAFBeQO/Hq//7pJJI8KMxRyj2STAiGZhpoUpN4cW51eZhdWLPzDwLu9m+Q8M
Tn0l2OrseSraCawRWlmbQMUxD+wP1wK04ejFEQfly0DjTEIm05pjHUHY3X8bLfgwHHuEHYSWHNik
SRi4WmrEfRcTU1C9lQb5zhwPzm6YP/++9fJtCtflqvJVrXFBu4o0tLMy2bcQKGEF89dFJKnr/HeE
WwViQPd4QRozxwzaivNOyqC4/rh0l+qHV8SWETZnl7F0njpcUAVkIx3Sk2OUFOUTk36qi6JdeP18
AXB6wdwOktksVh5OqHXW9vwy0OO+eSxbxofyBVWg+dRZ2hYTOa+QoKQZXjaV4K3MXICn0HZ3MwjG
EW7HxOeHFwLS07v4hTFsO9kFhpW5VrEpLEDMmUNflswaP4Ln9QKFxzDjHXlgsZZ+T0XUEtZEXVpI
VCy3khOvfy5QAJh4+OzK0oEF7nVkT8zovCY0oiMOoQjj/XokARtsX5TY59K6wtPOJHFKIedhKavv
WXREayeJPPaMjMRq0Czywsy0Fj3CWpseAzMB5rILvD7MxDB4IPD/EzQ5CGcAluZMFE3xvNdiJ4n6
zfbqCaP79TZpWtKAF39xhmSPX9Nw2OTfdzv+AH7Zkq+N3pRWx47QKEpOHR2t/2T7WNcK9xFkHa/g
23JOrR2lJYU4iAn6Ym1u5hb+vPJfI/OQUjrCmgEwRDFeRVBanMLTD6S57LOOnnzK0UQ/x4IFNqJi
WKGyZ4rW7N5f/tiBYeysgyoVQpuXTWbdqcqous0CH7E227xcZlSoS954/zM5SENEt8IfyD/sCRxH
e6es+g6xNg7ij88gPFMRn8j4tXQhR4ZXYVrbzrO3UtVc39tlwnjTIgQpqE4yDHuqLYzUpZBlvadg
X2YItJSauCYXY2jk14Egrw8aSASaYGlwIJyb3Xn8ndrGzJiy+ZUCyU5W1qUdtm2NWdiTcYSxCAR2
ionpE83zYJ3PF/tZSMNAxG+Us7E1Ct0ufAnUr8T7kw+EHC5w/TxZqd8aLJF2f6+XbS/C7hO+zlUi
LBgJPvsA5SPrSlFTfrw5DbWkVqthV6YIztg5GaS9ieCxaLRUN9orbQLq7rUCFzpVCYdeqW4n7tLu
tB8F+VJOSE3L9pT0KFls+fvKmRDoUAnIleHhcX5o95L8hJ69XPYvdmxsHyYf4L/adcIdXuCilsl/
DvGswuyfnFxCZgO98kC/pAry+PoaDcl9oVh3XmZglvdfCFy7qB8IBW2cLxY9lAYwSmGDM5Wdj0A0
KtiAnXsEhmS9fppoRoKWu2E/yFpjxxneY0l6ibuaaIIm00pQD9kT0a2VvbaK1InWSQUG3k2Sb3pK
Gwpvpo1q8f8e43Sqxzn0WPRyEIZ8kSi+Z7P5fXZTrjfDwIqYS64FQHrOVXdEU1XqSxScdEwMKnE6
zaLEJ6Fy1UHZDr3Nh9/hNeg8zLnC5/YunkGsZiUJjzOK/39nxFzVY/lw3L3jbAnpw6lnSpYifHPN
srMQetusMhLzmDLzfnYKTB7qUnPfZgqR+ItoJyOFconIMt5BZnbHC+3Ueoefpb4D5k642BnDhT1Q
4hI8xtO5VVltO/xX+XmTo+OqS58gEVleWPxaVTR4ZvZTMalFdLUS0Ki7uBeYXCNfX6K9b8KcPUcx
ZeUT2TpXjRnQywWMGBxIGhh34uHzXfkAE11u5fAFTTTJSjcLDhczxuYKthTM6qdcfw4yUg9znHDc
w7qaM84AeeiYIgnmRD1QPjPL5tDayxqQauZ6gGTkj6mKFAKNrDGgFp4FCmy4zUqPXd7icbRQMNbq
r5bZxmxmZ26veH3aGfav+RXcNSSQpmxB1RKgEqe1sp9pfnRt8FmrneqVvrQQUEJugVBfmWcXZMVx
J7DhTIvZ1Ebyvn1mAKaYsu7Jg6zm8oB67lZ4ehRBvIvmPu98oMcJkLFTYtXeZfHOQhyTW6+gSt0j
q672+iNgER6V+n55roY2ujKCnvjJ117rMDYbR1ozxi2ye/q07/jP5XQiKyTyhGrgxGwDHwQjWdOy
PzdkbwAs6mRhunpn1hgElPv/R+PKxJJPiF5yUi8K3smEXttQH7m7V3It6mso7K2eS3fTdlA8hg9B
oA1e0qo5I75VLBvO6efYIUWAkB/Jmz8hFh3PiDCb/B8cj8QEYJbcKAIgGpiKoLV2ly2vZ9qLhI06
jO3elIrmTC/OkvRSXOllbBNHwQTkQ7yYsP+y8Wzd4631WeclruWramnAQCZi7qKI+9xXvcg95EAO
BdqVGtHZ2uJUzcKM3Qco/LvNH+MdobOFXVsnEVvhvNtf/Bbw7221iX+US/QEeCxjim+K6/HgvdEC
AyrWRPWIoFMkk3w8iWrVQpiwAXaNv+y/Xa/Y/cI44u1vhKzTLmbRZBz6xNIqX/1Dv0pxENIIS7pe
NHeSeU5uBxfZKHNAGBXppZplhus7dy6EuZB0F5omQj9sIkzPKxWyTGBcgliW4KEmGadKKDMY/MsQ
2p3WdN5SfN6aiUz83H6xJe9lwMyZ5QyOf3gsw2x3O3VPPS0BN2BhlJomWARw3I7+ukLuppsuLB2z
PFb6EM59ND6XwNHMOeiV8sDp533MTd6a1AFIa1i8jYCOKjpxnjTPssLEVa+i80OSZrKRul09Yfz3
++TQ5Dc0sA4tb+z7O1JiD33LG3HqHTGcee5g+zCY8rXOpOr0IejIiNDgSZORKRPGXEXGtCN+t8bG
lPjAkAm/ZoGm+V4UzErBIDOV4vFZ1ACxCN9eMf8u8V3gCtUJsgbzCgOOURd8jNpyCsSC2PxVqEJa
lEKDocYfgAENqIgDVhgykQi8noGiodvPg5rv8xhdV5lwbMKA3/ENLbFYQl85s9paWF4/Q2CFu5z9
RcUaxiXBPmEfciEf7ZzWnOphd8eK1BSuvwUcpz9vEWtXYALoJ1tGY0h+El12bLPVr0L7fkKGnucr
AuC+XHHPNwV8F74//LVRNdZfFEqInDVeDGNFMdhgpXrEASQ7V80noXM3XwuSbOAow+7MYn0UbvAX
XOD7CqKFpQc8BTG0d5nTwUloDYekqCctgxenKo1ri1SdO+WnGg6XV5KwP0wBg3c5YnByBu9OaQ/1
KWhleibYjx4NoghNEc4yOganUUkwJWcrhiodwx1CYPe1s2Jn7ljmnVA5yQpchft/RdZ8WJPymt1w
NuzqfsKAZVX5mP7I5bxKVONK3c/eanjl1FjRt/xVzTnP+dKKmCynZXEji/3bOkLiGb8c7wVbrIlW
adiHCVQmxbX0HzmGUSnm0tJkhkL9WytQ4GGq3LOS9JKlV2+3ubytoxylpxv7oP3QOiXTcb7JZNLx
P1Unyed1lAs1GJNzvZzHu4cpNTBoQw1EfMfATkmF/vCkYjjYrGT4jp8o6eUtgXEUnXNNK0f7hwqr
aCYb7pOH6PiYbRy6HwUpGo1kEpHDlUejcBIzNdbIP6euBg1KKvN6wSNB79sHXVUjnnls3BeVZvYL
YczEBablFuOpELlgknq5oREnM5uMp1/zx/+imaIe1UjxWUF2ELgC24DqbwVeIvu+g0Uip5/M4CY6
vbAj8sK6L5BqBPHRa0vVjBYAWS9ORhjWpLfUddGCSAluhODw2GPGGzoojX441B4yoX35y83lXr8+
mxQtUoWTaLADH+S7wsvkprhd52VgQMCu1NXqMIeiAz9GC2Q8wzLZgxGdRilJROdyeb7hpD76T6LQ
rYBsW7IX8vmg3ueBSUQVoUFKe91HdSzjKxBgUpLu5DByqWT2tnLtAduXBufS6MF6J5GDvlNTD4EP
lwdjlVL/wzyw874jU9evz+UZyMHobTIzifoZoJi+rW739dzuJIwKAmGO3+8ehy9Ua8oog1b+P9po
WGttHY7XDXD16Z2BvKO5ApJkbFANN3yLQ8CKMYj0MseblEXpmYz0QhVt/hT0Zgm4He1ThQtv2f/x
tiU1+DOiOINOwUslmlMVq7ldIC6ryWZgpFXvQHOxvy+8aXKCTa9aGIdu6fz8U0j6LatXZKJVqxDG
kOdXg5YJ2Iid/8W3ngV8c27q5lX+1I72Fat2MW+PhkCWl0e3xpnjM38nX8+gNp6BUMY0tJ8bpyQs
xbNsZh0bv+N/W1khZ/BJ4PgS89i0J6lFZT3NULdzCo0EyiayqCKfg/KmuzbHr4t4eEAjntiL/GWY
90IXwJhsFPZ+BuMGiC0035HY23wE/F247Zmim3dxDmwEs/Aj5ilvGwnHWwoxtaYTmZ/EtkodmTjb
1X6bMegMT1TX+hcaD0LOU0MPa1k8Vm28taF7+HjlNMaDNcglHoaHkcAOuRpyo7zixx7We5mkVldC
2gAAl5Q63NmqmItIe0JCZssTA/SwRfJBqGGfvW+wAt4qwR4puxxOSLcQsH0H4dRN4/OuwSUoYxw4
GLcEeZ9w2lG5K9us6PpS41ag0Mdvbycjc5be6QvJJt2Pl32yKGFMIUiO/GeeLj7YcFqmB2hKnS7p
gy6CtKAzvmreLk1yb6cbRNDpo4qfAL45k09zVmWPkPBjEz9K6Uuu+s2CiEUrbswjtjins6vJSd9v
5znBecl5lUjnGkbtGJeubp3dG1nbedpes7z+HO+5WXOHdcCo8b5NG4a/0lynmDlKpGGJ1h9AXt/d
g9FFGUZnn0eSmlIkSjZs3j9Q/38uS8W4b8Yv+yTxqqxuXLuFH2up78Xbjed2UNTSSjm+r7gXfZ3T
bHNIuo0ZFWhynaAEZifhOwlAHHgHiCkT9Q6tFuDGA4zNWlNjfZHNboSnUrJ5ZjESXiCSv0axYJ+j
miCpeeN5b2+ppyaOXhpObRiMqybZ85FyhUKleomPXEq5HK0kZKzt2QQknEf56P/iZXhsqzZhkuOG
ENE1vqg6BZWhm5jF1wKJEK5t3GPIMdLBYZUQ46h47zcg8Ppo9NiTSP8MliFB8QLaTehxa5hAjp01
kd8GLTScVZENZM1sWw7jslwdSKbP/tPpZyLMAJfYhjUKgxf4N3nobXUL8BLTK79vqe4RVfOmzLCg
spDZwD4hpxfoIFS6SXw28e1EPEZ+XzcX6pT0EAIsefpRPCu/SoNcfpm8K/1S1wEtyun5AfHKLR5+
znpPOWX6Jk1AMDdVce2pvJlq+awRl39YZ6XkBBSZ33EaBO5AW4LFNCfQKG3SM552huXuqX3X8ly5
Fv9ZdFl+X42hgJcE67NQcgMEVGD7L70+VJif0X7V6afwGnd7HFHwCQx3h//sfO76O8V7F3LNRGQL
g95A5VHqx/Oan37s5iLLKmZk7TGT0fU+h4ZKVPJDVt20cqBacjgNkF+jtr1QBEpn4IpXEIOr1Vfz
2BMngJshWg3vUg3tX/vd9PL8ogQqWHem8UlM2lvovO/TWPCfr5dzpOl/le4Lcio0bLZkdKar+I43
bCuRIIr29Zs1woSgSk6leSAh2WNae9aNULXkDNtQEIB9xdMiFiPWNpqauWGhJiXs4sQ7pfpX156G
Ldw8kGL+9SndIjr7u7tolzRaFLGjcipKdSKmAZAqROZbYcivKv4Sk3POMMefmdKh9rbC3ixew1fa
DgprP4YXMagcuj+DyAmWpI2krlI5QmjGefokHONM9tvrdTTtv/RBTokQ9n8J3c90gdFoSaF6FbhM
Dm9f3ncpadSQCZxHtzNJrKofnyO2EPpQRek3Rl4Ve6UfUIgv+VY6U4d8GxOBtw/sFgvffDz7ht3n
6I4fu0ibu52ZP1aNja26tBB5mCkWnQjYY3LHcs1pMIvfRA+18gcA9OMrR+6FtoKKjwRom899KmX2
RVFYFkkLV0mNKYqAeDlPZz+6hG5p6dHHnSzIHpr2dKCSI66ctJxGPjTSpN2t9dpfE0fqNqO3b7E7
YHg1yarUGPO2DNzkesy9kc156MsWvWnRPNe2Cl1eEozNS2Og/ev8ndYOPCchzc9rI8pveIqNJw+9
XuMIjGLwYZvVKzIZJ5e5FG8M1y6ZkHwh2Lt6MHJzlc10LrHghvwaV5e6bhgZCd4bQ8LlWXYjSY4n
HLkj9+RGhz3AQq/Ar7cxZX4Z8B7mq4G6NdFzZF/kDjzHZ52sEtxpXoewt++Af+7/XeCpw4NiT31D
dHp1zdTe6bcMvgT2V5EDTcJxEi4ExfzQm8e7Q/wAU7rWWuTjXkuM0iDZ1L6jl7EC1wvc9zWAz+0j
k1KPQbvqln/GOwuihicBmZwQxsP8sAFCr0VVBmQxvybUmvNB7z/gQfyJwPgJ1HWoCGGdRhjSE8VH
7ZUf45Hr3Ad3iHLU2cv80l8s5F8ygQFhhBDE8aPcPIX54VE7Isp9cJ0JEA+yfD38xwIWL3EW6w2w
JnCpc2K4BsC6T4daiN9Frm/9Pywq16XlUBZO65VF0/VEIM4vdBlaL7gNFMPlCSN79gDKbIy+U67D
36S4LkEA8NuxOKpoVdhuFAm8osyfExmvCOeJBpXh2fkW10hMoaqLFlEYzQ90XsE1zgDWnsUQ/u1c
fGpZraQqo+/KfQc7My0w9E+CUBjlTcwTYik8WWrVZLza6rdrJPZwDRjHfGy9gyycOyNij2uRj0nf
Ed8RmI9adkRa+UhARH25CaFc+t37d4goxOBeD2ErClb5LzvWKzWAHlldXajX6q1El4UltNNVf/wm
/zihvbbyjzkNf6qCo/4SXJwwWTkQRSrAbqnO/s6TeJ3e1XSzNU3sjqGCco6BDp8U1MK6HV9vZu28
DVyP401ZeNNunQTZymF30iQOlGBl5Wn+h1MvhazyPepSK1qlvxXABcp/M23/Tamdv//yWZcwV4Ix
+5wbLLndI2VmYra6W6PWHkfi53N0a6LHcKFwSoQtnukLGoE8pRt31HYLVlblLZMrU7oIZdylzMmP
ZTCLKH2jl6S0vGkEBBww6iLyx2ilYTm8Fw68rBY947pp3klBUsiYKKrkIgEPHcvK0dqPWMkptZ6L
4vTy2cM8yHmMq3lKPjLEayjVmzL4WSMpeFhtAKA4Pzzt9UxMWSy1xvDgKIVboyx4pO5L8YpOLK7h
LVnXAp4Q3+qx4AVwqiXOKTedmQtm5O1nMmWiu5jzgDhZuQbvPhQ3cWuYoou9vQl1cd+j2Z3JtXEH
yfDpl4Vv/jDsEc5PvdKADnTCpjpdtJvNmJeZycEtWn/5IdqIdudtBFqNrGJj8LR45P+G0aJd68S6
h8Bpq9TPg7ix0y1Cy2S/oR06I3jdW5MY+tZR3TDK87o7p5gZmlK4fW4Hu58Sm9dnZYBWFvR32CUZ
ZkCxos2tcuL+vq+e3h+lACbEFkYMp4oBwKxwM8UeGTI/RDDsmLwSY+a9RhwYqeZIaoidXWZsbkXb
/N+IQENhL4uMw7cKKUlxuZumEIv0xNp6eS+d4tE6p3xHKLtpSFxhj1T02dbHxAlXqHzBgcC5/7FC
QLEvnQkqFRpphKEwdp7ZhebgLVQfe5KRbGvZnLc7SorXRVvbo4M5UzYudlxZjTbctFWVYBvyPhb8
IN0CZPfbzsRpeHct2JwpxMv/Ck0u28xEXL0A4/sKiIN3ipfoH7t/Czw2Pvtq/gswCdBtIkFpj8t5
FZR31IKziHyFRL2obBIpTxHNISImJJemBtjmvkhd9xx0V3cdcL3cTiVnwHQw4rBwvTP1ukadpMGO
x+U+6PLMqyqrHVXRWO30yeXeyHWZaXrVO6/Zw9oDjSPi6ri+3Nbzgu3/ZAGv4x4ZiGmxASJHQLRe
qH/9ZNsbuTO3WB6g7o0I0g4Z4APx01X2665UNGsW2USrFJfEubAc8yl2MmZmRpiKoDJMlrAxOA9L
OOTQ9euCzgPWtngL6u8hBZ43F8+exZ7SKOzz9mRcrqztYrwlScmw7WJx8j/jMGYgXUBve+F5FbTA
JEPN55uTEq+xjJitgkUP3lvBqkuH8qSGsc7CuqYlCt9xOgxFLyqU12X0nAD6VbX+cba3d1v0CHn1
6wT7i1WO9Sk+lO7xAKMmBC+xMuSJTdb8MHASXAhtDyRnZB+G6fxCA5GIgzsjs17OwFwXGT4MqA3N
d30xEvMc0lgu+oHdpab/3h+i28zWeqg6MfDwXf4HADb/xGTSgzITVdz8poSCrRqQIKnHigQlZljF
y3m8jUW0NASwOLG0R70b8QFIoHySzfkyofsm+UDuGuCjpVDW+kGcsXFdt6KM5c/k3Y1KxcEixt0G
YbDzdZU4ZCqDzLhxpx6r8yJ0HgYUA+yCBJpsyskFJhdjZHLjybnbXKwfHGMK5x4oX+RDz4agUeeE
eP77lnm8EgN4AEK20grbHhYffFaDQAy1JIA/W1dDbcW6kb7P1iXAQWs23gf0E8jE8TQSPavjaIPq
1oc79Orynn+VtqUincGTBTnBWn3LtbxD628zMukgV5Bvijq4HBYeoDwPEChqmCE8rSGIAYPvwHju
gD7Ol3lrTebP23p80DclILyfFsgfFLF++ZuJclqft+meV4a6vkjIlZXuNEd+9+QSLxLoUvdBQdYU
0mimqoBZXsHZE790sv7iYpFV/vvuOEJ+8QjFsPFpXOdU1rBkPgO5yRZUQgMCsRjvIJRLZaucvR58
DNHg7lJ9KM5DVTlLU4IoAPdJQEd0sslZYx2w3Gx5IVgtb6UEQPBBkoD1Ta9rGT0/wEBcArqlk9r3
bOq/UYHSyT+WW4aYrJMHf58Z6gDMjxO9F6MHoCxb4n7IsrJLJGK1O7vm3uIZKQ99CVyQ6fourGg/
bNoQtEjtHab7L75X+KJ71hG9CbHbMw+yTTY8WxF64ttkVgadd75TytUOkQp60ea1zNgFInFXsyxw
yFXtbagrfVFo3q2xJWtX2EiDRDxy01gToQOdMNUIBZ4iCdp2c7r2VvKy7jL4DYtWQK7exRlb/rQJ
6JK2GB9AkOlM27btev+pgERjiIvnkEUTbaJInLsYoGAfKIQnm+1Zf5u4YWPSRrUz4jcC73KG7aRa
hs4kxTLjoJYBhLndNx5oseGWUC5NakN/P1SCXyQKX+rCJhbWG2iQBGCHCQHSbL9L1EKxVpWoZHHA
5TLsPC9b1ir2k+MNY2RUKVPKxURwt6pcYK3dPQEptBYhwdpuyfi0anuNiyodWZybjYeU4XYtNGwI
0OfjIQ1E8gSS9RbkmA1BNPcBUoHpioktsLxmxe5hL7r1mnLa/t/rTQg0OKzPdvLq4Rhxh1498m1X
R/zxrHgF6KPOSKS3+mTNAIK/ThIDPnG5y8R9TB9AE9Yq7R92RYI6GpKboGEykA8qPcpjUJr3Ur+4
AhXHSLz3mKLenL3iDdOFJe1dQKU0SDoEsyWgQf0bsFNwriW1filhQ1zP9wkv6QTDo9gUlDZGI8uL
fdR29XWovbRD/E1Zo40GgzQYLX0kn7scQ74b7vVF3W2DHeJSuCf63HnoUhOrw6NgGk6TOLd8sUFZ
zkPmrph2XI0Z8eV25srmX0q0MKm67EWmyLvHkz17AXT4NQXaNL7Jaym4EwPtiKljLiT5PjYppx71
+idTaOHkO3Q0Zpw/tJiUEucpyw+mbL5kXEkpyQol3PGrKgjslSn4FimvHqf+5T5OOZBtJpKjXEWa
HI9rnI+BFXtsCKZzW1lW4I8O1l/e6mMLUEahEJ0LniwrnJXHf0s0bcypP/dD3qg9IX91m3ZAK1Bh
D2sLLBvGnccN+qCXwm26DuxLh4XwfZvkeAsSweHcod9ern22Xu7FRrQK3YnNPH7vnXmEEKItk+oM
unsHnorono2GCwZAHbayufmDLZG3+K5vv7W8IBdTiFoeoh1/m14P6n2WoZTmqZAL4ldgT0h6LfTn
m/eX5G9bnATcoi0srZtLpOgp2e2zId6Z6NSkZADaZ79hXSso3o4gFjMzyHzgF6PivDXkL9Gs9rfq
JCepgCEtVGwrCjRwkjyVuSvKPxV0KjiPJx5p+OW6CPU7L7g99wkbxuNoQWWa11MtngOLx5XLkGHB
z2yAwCB8v8AC8T91YY8Y+kITfhvnWoXe4eHWmtXi/kFpJbBi2ElUwLbhp542+uZ/vnw3GZjIgFr0
dT41q/y+bapLuzEZ9B5fx8R+se0nIMVrOvvhTtFmdZvXaZf+Adb41zsTr+/9sPXqQKyclPnASYt/
ruZBYXZnQaKFuKXmJ5HKUaYSJbbvmmmgHIImA7ZWPON2wdy/Pezp3GRHgNhQtfPs0F22JR5TKoSd
juNlkLKWFW/y7VyzsaYYCkThjZnU6WY91IGwFavEI3FwjOYmymQkJIM/FX8ydOvr1CiXCB2rDGG/
Lc9ksyPy0EAYaThvdREn4D7lDYc5NkZ2iK6K3aRhNHEe/X5ddlhVljcvrAfhDsiF5tMzrA6q1qjP
xYJyIfmy00gFeVeGgRgfkgwoHjz64OJAEkH+XTz+7kNCNZSAPSC8IdGe4uME9V3H77MNW2Hzxfxq
Rr+M4yAF8MpIQxPfoIecQRE2ryphGHWo41owLAv3YmYicr7OZk4mQ1OAcMqXLMY2hxJOpueVGWvA
DY/NsFjBcPHEdR2X3gmEVNMiPF2WKgvCGKd6huO0vMiG8snphZlrBVpa8L3ZDpCD01Rz3Aaq/+6m
3SLCqKz8NBRivVSrP7UqVTA8c+JQYwWA7dwMQTTFHhDAA6KPBL0t86YTFhAKXJB5PK6U38QseQ4p
nEp68t7lYoMd0CvYE5OCUi9E9xKIK+SO9p+/+j0YRT5i5N/hypc6977dA3s6J50ZYDL0+8fTK2it
N9x2iyN4QhREZw6vuIBbSBSBBJfkVxf1Y6dswG8+0eIckB4awhmE9yU4os1uCE0023SdIbPGlIs8
7ptVoR+J4zsdhjsdpm6wtwdw0X3NSdCnjcrLmu6MuvgJsN1G4xQhnxGIMS0qtoBQxqiD79DyZ7F5
jHRfB9hrM8QlxcM4tV3yexh7nsWhcB2wsjswiMqCCTQ/TKfKaFFRFzqZf7sPMSbTFlgGh0aU+5ot
BwqtCpg/+F174h4ugASdvQxYq9+LSgypE6YOFu6hC07LlQVgN7pkeDozM06T9aTg8xBBawaKC7tU
BFPOAowd+XyqhPin2UUrV2dxtdLbVulKmjZhY4UGol4gUdbTJjd8X+fbA6hV4UVWYXlaOhu+WnJk
/aqy8+0BXSzx10dqofHz6AeYJWrY4EFV2rCyQz2gqRgUdFBgMxwgC4AtIiH1FCArM9XJxwSERilg
DKXekjXgEcEuLA7OjxcPj8noPibiGQFJP6VazYZnfNGB8pm/GIVOrR95R5lAIgXbO1eRiItl8j3z
SKycGRPMny5TNP2kgrkLKTkFg84CAit4Hwolc38S+3EVTQid+BGm6OJ9fP9mIB1iD8gMCuJ8TsiX
KKFLFYeEyJdZ6t4g6HuqgRk3iPN20dtcD7JwJnA95FNiglFY3zy6Mn8qo/TqQRtks1iCW8s9DG8u
ImRG2r5AR+BdOCWTtJb7BGzrCebdTJUsVWvZu+FzNqwEZ5TTfT2D1i2dY8sSAbStfePLeRXKZU3j
wCb0nyyPJ70zo2EabK4OlRs89CxWoMer7mlwWWgvAzmXjWvhlLgc3q9Hj4/sHuaOTP83nYxLMhnj
2LwJo2CPS4lh+SMLyhji3d8YmjFxONuI+L37cUVwgpzurWa0qt2RkernDzrJUWTdOwkeTAjykEWF
L3/XJCPIj5SCco8QC2+eP25edDy2Tn1cy1SENR/QxT8r/8Cv2R2Th5rZW9zrc7CzVigjGUsxKGlB
O3T2m2EeImyhVIR4pDb01CSt1QQklfcyjEFcFr40wtAxXJ+BoDgFfymyAYi79wXZu9aQxWQhcXaD
C7ghQoK+ApIBaPfzx1UDiQzY5Z53XwwrA4dLzirOYHpqiW5MiY1SSm5nbQLShTdKF64dQdhcvPOO
YfxSdYnxZ4KYHU3symy1Ds0BmaC8XKrCbToixp2QOaTRN4gTGc+jN/+3naeXT1qdIXJKfM5OmYob
dk1JCzprYEbSqiosnQdL5BWp8sSeoNGmp4dbs8u8uKwanhRZLOSmasg5AZ+FDiQCT59tHrIYdf1r
5yC+RNlh3wzAvmfM+WcxpNV6MNGH+W8gi4HJLB5OouJC3vjLDZ0nvKmZghaVzGQjibztCIo+Gj/i
XZbeulA+tvomG4kT6TJNzRgmx4lBCU/usKWvoAj6K6ilN8Z9rpDF7tHO8XhM8mb8F4Nf7il4yZLL
NlcFc99kFwVP592ld/bIUkncyaoKO8CgMYG97YGVJ2FzgDC0anP51fGRrHHRmZRfVgBhrBjYU97u
fDIkTw9uljI2HpAW//KfaUPcYiQq5Z0ChfwTIkR+HKaolbeQcEanSce15dFRGyMUvaM+Kzj4DtFE
CwOmGaMSIn330gmBpT+pMToEmzIxE+Im9mZrVNelrRGpAPJZ0x/isFh3vaBHIKL2nUMCiTCnFUGT
2MoitVh+RhTDWwi0LJhpOMDPR4Ho12n+u1AS1zT9eknWx2SwIZ5icYgMkVtz9mxSIAFj8OHdyYeb
qgLWl80J2pzCF/dtSCBLuqp4CMu7FYr4YNzWjezT3/DEhuev5JEysMhOgZlBsV5iwf1nbNPm9bfu
MtMjGyOebNVobk8asTK1dutxpt/mGs04DTCNSHNKVX2ESCc+oa3COPHn9PYlxfoWIvfvYC9+QVqj
NAMi26d69u8mwhkviTMjsnSoOSgd+lnCnLPyOPrQdNTprt9sIIJ835YyFqvEfnVD2bmasRzQDhpM
pSS/3rV4I//EF9Msw9d90YNStMpLIR5HHvxgXpuuMjMhDxJcKVJo6wweJ9Zedv0HZoTzgLE1AOno
a03DkYGTv2sE2OrY9TmIwjMJR2yMM5xgZkIHQOJDhaHOfBURLBU9FOj7+yKkteuiZA7Lqig/qXOj
m01rCiWABxwsFsYmLNFGcwryNTRpKKGNYb1sIbBzZR7zply4IMZnDVvEGkQjMP0nZThKM9QeF+xX
g37UlXi5bPAMPc9sfK23gbRC9zbZxVGFPj/ohSSkXkesopUgmn8140mcimBU0qsC4uQDGqaANnMA
HEfd/gwC2gXgNETK87n7NB6prFBdNawbSvc8SVJWIPmq7JZMNgbvIgxnK9e39ysbGihPGQ1Pfztp
0fs+F6yFVrsdY8ffXM4GEsmGEYyNdTIE4Gx3blKfY9pHwVE+TcuHdeq+EUkjMLPsTTK+NQfTRFF6
mnMyaqLqMXWSj5CvNkpy1km9H+7jUzzt50emXd97FiyEAOOGHRBp01cv1TRvWguz5SNogpVNnu94
vgRV5uMvK0vMz/cwwcuFimxgaSlkEG0Vnq2xOoyofb5jrZVW+GCY/xIoXyqrozlEDs+o9hMetsKz
7T7JHqH9nOKt4TDhup414SqO5EP7rJNwrCVhtV3b4jRjwb4mqHEgG/1Aq8L5NHzkfHvaxQnFRkB1
PiVugMBCDRLAcXZj0PL7wUX1i9OIyTCIstUTK0yPGFkSz8f8LCHocaU+POrhgQhKpHTUbkejCmdM
jpHl/d/auVKiQ4pY7CfPVB53oVTuu7Y3qZfDqmW1kXj4i9a+yibHaX6yQc2+a2HkTLgj/WDwT7SG
ALKCo+TMmVb3/za4eWRDvbJMZlTNopLRZuTqY+i7G4p0A37A6BylE0tVlaJIhpu16yFYdTJEwCC6
Vp52FUxlaW1NeqrmhDasjwwbK34w/CF3dWXt32ZJ7LJbnIbwRgsreYjmOojWCAlharp+8EijS1jx
sVklAVk5IXLWjeDZ9XszJvmBYeWmcHA3ujOZv++ONvPRsTbsUkbGlucWN7nEA3NES+TwYJpsX0sY
TIkicW9iJ4+8P2lBZeg3VKbKP00s0PWtPYhuP/V4hSNPDA8e+FWLiE/acCAewHTqQftDfu8nlheK
6ncSrMUBf5k+PBPhUPRHRAmQ5LhgJHIZOuZepRN+aiTjqs1NglPtAXBvouCxXITnNdTqsiLh4znN
czMrGwp9TDh0iiwIYoNUbJEtx1ZQt0VuPm147HsfSyNmiOUu7YiEbVXVYxgq//5c+zIND/NBdTTl
fn96NJ9cdhluLcCp32xTj7pOwqMZTfKc5MRT0WAs2KZI0vSkWNuoKmZaOX2eVFw15o7ZbfB3eqfY
PAvnHogQL7+Rl+26R+nNlJB47ufKIGFQIWkmYBAZ6Lgwp5wdc3N6KIRuDxajZ/u8KJAftVjNqwdA
q3Pd8fXu7ngFfyGvkgz6x4QsVTmB4kOgOGUARwHbC23GFUxxg1nFfxECWUY2KJWZe4dX0iJMdh9O
7/FSaq5E214GRYzjv0e/jkrYpn/60qfcOlXn3/C6FsOvH9GTrzTQniErxzwBiWf2yG3CFBuZ5lEC
mnvGeKXaXeRk/yUXHGwGJ8RrwYz/kficX/kMdg2U7b9uJvP2ijIEebgIEWG2to1udrWQEa+92kDu
ND4sGRPA4QPvNmYFvHAA0hSbshSu3teAp6mJTOlWskcJmlhCh5i5kE6LZNGzxrSKw8D750FJccfQ
HIV64IySkJlSkWukJgWIk1ZsoBgNOXcf8PuX33NbPYubErbBtLqOfie80idDc9YAr9rOg8G60/Uh
DyBCvP+4mMhT/8Tt11uSLPfnGYbZd6OubE+icWqGAd0CvLV5AVC8flh1DhiJuI3X+v6h61+PHUol
Hz4jF5byZybbnRZEMkGZuhL87gf58ZL3hHX/tJa+++QwlTsWXu1Mhr/oVmDPiAPm0lappi9NA/cX
NvBDrVaX/7WSFC8GxVe1ncYK6YANP0XXxNG6t3J7PyCFkpJ++Ciu6FrXZpblulWCTXcoAXYR4dzs
lzq8PFO67nDNO2GJ42vz1S5oqiZK2U12mQulb2IfnccraTJxI9dj1Nzeb8CcC/oL/8xuz+yZcG7X
e3eilbwjMIcLxD6ps0SsugS+CGjdymn6ly2pYZc2D1En0QxlhXedQuxy7cABPAT074JjubPxgiH+
tOhbzCoML+STdo5oy4ifcBrPja1W5SEc2h8ffHfo+yNR8VMXvwAgzaFcqkZcWt8BiCIL6uacGUnz
ZXhoI21hPa0JwhE8ZS4h5q/uWWCXiHaSd0uSdj2ml4i9D3i4nhsJ87fEB6wutXh1BfzYTxhElumx
vRViwTmKqyM5PQxHBvFMpBGbdjl3cUevbjYkMZNycA/OnihLSTkR1O4iRTaxB9z+acNXFyH7aH7W
4KS2tYZQUVkUk910uN7X6u2achIKrbrhGwTIntRaEnoSVux1+QrEHszbXIDQktl1emcHEGDWPjeC
3pcESerKGPw+CCAYskjFUcFI5KIEnilndPywXGqT7vZdFHOs0swoaV2rGZfRhUNe20x8FBhMAJHR
/TD/UBkNZm2kIWymUnOK/fAzGnx2izwYhovZiw+ysLiM88D2wvahd3rLIkDA89Sx1L4U7mNANLeb
+MjEm0aJfEjAShmK7wD2c3x24WOYs3A85HwD4958e5uTQMLcp79zFjH5mZNPHI72tiOneouMXBiv
6LdbHDAkSrM+OOSjl3970AkGepyIKqx2gURRBQq4kJj/JoLSw85TO1Cm/h4MC9fsB+0mx49wC4jP
4MdotiovtXxrc/jtpsixfcz5iDBuNOiQGdiD3HT9+jV8GH9O/GGTKJIPds5o1pOp+U/qSq9gj56k
xVYZE4A0Bj6JZNyCOSUTWLN0uOHvqiR+Fwaqalu2QdEusA1pfjxPzRUaOk0VrnpVaftT9Oho+frf
124YEnveKPKvC+YSwjjXiISLzq1VkERulqd78/W70x91Gr7hpelvId/xh/s3iS7ZlGcJ+y1NDzee
cYTQmLSxWSh5WUQG/oG5gMC2Q8fUr8fJIE6h0JfMFUglbAkWE4b6xyB6dpYYL1EeOIvy2heQxG+t
3MoSvIyx7GxWmeJZWP+ZuISCjzhSs9K/xz89MeTcLXnbgDpgmNrpZF5uR8dz6FGnYlWJIT0WWX7c
4+Zxa9QKfLrM6VFsAvz0opxjnxoz7HSEIRCRE30BBMA/mtVRMDneh9kN54UhfGpt/FLHm5NAP4az
ck5IwD+xkMTc8MWup8mWkE9yebM/aVYK+JobyWR7VI+F2Eis/gu9lJyN8ZDKHk6FJw1xBbYFR5oT
NGXKnZ7KQr1iCIsECf0fZvgIiW5y5faQYI+BJSaYqMLhZN5uy92N8j9sr5RFp91fdNDgK0mUlaC2
bZJ8Gs8ieHo0nJceULc8YMOy7ETe2zjHVhuqR49nSyChTCuJmKNEAtHcCxr5TdHSn5gMv7TBvNMi
o+u3iW+fI4enY1S8sjtM9XGi6HyTdeR7ouxbGuaESY79aCrd7O0tWRaB6c+PcusfS3ETTISL0O/0
/+Fd2JJoE+MF3GFq84j6UCCiC7+malc44UMLtj2Fh5Xen+jm0lUfZQ0w3c7YeHjNdu7mD29XEH54
X7ADUeshEnZvX24mj9LvpHXgKK/mqWZTu7j1EEJsIJKaXxAstzmI/Jy3S6qCPIE31Nr3WnLluwYT
hJmH3ym2yM5YiJnqD6d1FRoPy/N2nIRbdnJS0E+KMt/I6EoUJfPo+1jLIsNEoz96pLGQYBWB8nRP
QZpIQ3UVGRw/1lytHKpqaSX2C4J/2YBOcb0IiYy/GIkLTe8u/xjbqrlDWEm3j8DHBb9LnJ3G4aL0
MXZBxE4LWiXqqtQJY5kYWZDywKxobF39Ah67rK91ls6ncXAXWnfFEqRzxTCUT0dU0RABdYkWubzr
X2EaarcanCf6LFJcTd4xsSplJwzdQtMC1pQxvyG64HT+Rh2urLm2Tq6nvt8Z4d1v6AwM9ZQH9DPn
sQPFmXCrORzWnI7ODEPLMxJxZ8w6VetRpzNIbJ4t1yB1y0xvzs/XtVyr7SdRA1IqPF+OIqy/ocs3
uVev87wslV7+9K7Pwri3l/ryDvpP1we+80e7qPi37iNErGd7HK3fZlunEZI3aFN6ZUiTJdbmsPEL
unyC9rtYB9HSsAXcFmIwJ3WUBjtllU77oqgTckXWPHwBzVxOkc/91+XRXhvzC1gJE1hHzwZCGoH8
pWJ+IfB3ASsIfET06qk+N0i/jOdxYUju42X33N2aJ8A0zJaNkCN6JX/P7P440nwaKxTZuFb9P0lk
b3jkI12yprv8IiiBC0ypVS5A7BaKecAAgKVcmhXe719BOYVlQb+4qjBn0lvfKMoDFHh97PNZn64C
96QGUZMHImxxQzCSbLD85ZsQkJrbOvY5A8ypHaJPjLSoWSjQs2tGZYk94QSLcITMJwCLGUmPfGyi
VRIEFueTiGGirrJkHM4Sl1QRimXtdU8K9K7hheR9lud85+9V9lzGw4vKIyCgl1AlfQPNUU6vb7xZ
2rixDSwhxjbdgarv7WXBzoKB/Zx2P3Tm5g53g8JXVDMORWWcuc2m9ZnRGOqQF6xc6ZQu7l68qIry
BUGbzUS13oJrZJnF8AREUrLtA1pMsLL0Gm+GJPetXD4rR4hbnsG7La0E9ufLKucN/C/FjBaASHPj
QICTy9IYCvu/8XEk0ov9TxCBAa+ywdUcZ8/4hZYuRn2QgTjoWs+aavJKTcqABi96TN/egyyqHJ7M
0SUbSUGxI23oxxPnp3PR4xRGRcjgbfdZtP/Tj0Pp+oT5Mvs1zQoJVDP1Uk7Fm8WIUq+Fo5b4NAz0
BsSlIkU8jz8dPTgGCq7hKm434+Rk9kipx/CNLlEPAHCEOwlVelINwkQGR6bObURFbIy9f/Hb5jZf
+3AkjN2g3MtOrvKjh6mrUe5UU9TQuiWx2FmmYyGrARTk4a0Ld3fw/rOw6zgSsZzP9GIMq4SkVWKW
tulAS1Ryomf3Zx437Hn6oWKNLWZ+seF2Rva1qIMspNDmLUQVEDYA6dCB19DfyJY/HyRE8OqYMiZO
XSxsl/L8Jj5pU8pFzYRV8JQsKtfodh1bwyugugUCTb3qU8pzanGOKm/Zmz9Ho9GYSYYnjWu3IFtk
cDwlM8YXGp9mxxz20T313gMeft4W9Xrrq94Tj5K8adQ4J+dvBvCY9W/Wu3N6sXIYHt8Dks5ghRwa
86e82gREaANZuZTuIniBt1q2K7eVnCC9jz6dSyuGYjm7ZHAFnx3XK5InWIqGmhymaLtvq7ZY5st0
nVeqJ6najO86gXVoFCcjIfsEod/pLBkYiiW4IF2Cv7i3+8Yu7YsNeyFj8gScpxwr6xqBvC/Euy2W
Bmnwxfs59qppf95+yIOjpyv2olMDwSoyO/Zy/pPT9w921R6pWSzXDPRBVO/DkVvARgmQVOQ2wNW1
OZsSFSV/E4lQNeDVAeNeutGDLWr9tWkvGdmZ6vpr7QfOIyUNOfFPfcyhBlvDTs8aT0lbhf6cD8Ot
X2/78MViV6jojwX45lNtBHBlDJmA26S5y3RJK0yPNo7BYx3bt9f2tWgCN1i/WgoUO0n9Uf1MAZPU
Yrw/Vg5IsuMwzCmbrL7eaLFX8M5VOidGz+8A0qwckldh4y8Y5ZQeFnLSSlUC5Eg76APEx43ZQzwu
Dw1SRLEhnY3dHonJ75wk/eEoL5pGF8paHuXFQuem52KhjjXvP3Qx/QiHPO2px0aTRAh1ePjNXybe
klIx5i4KuTwu/45Ex/h3lpNMjEdCS00ztryIB+9EJRbbKjJyohGq6QZnZ78sG1m8VxYsUYsM6nIs
Pw/UMN0EkYitpcS5l2zXOvTXnwvMTEdv8ukJ8wFZ3MUqr7ftsVi0VcOq7gy+WUTGh/jAidMnUeRJ
0G8nlJ00GHKA8ScufFtIe7ozWv1Fb3qV74NsjUa9eEuiyvnKMGeq4fivTm46/xeUxgE2RAOxqmb3
79kuTgYgqWKmV3Ci14C7WkcZMkzaIq1WhW8AjThnHwU1MKWdaJR8iSjxD478a1fKr2lxTLgxFMVB
8220y8QA41a0OTHrcof9arvwM2BZFdqz0VaCdiqH9N0zf/ZbjzTuTY0Ma1ivnpEdyasvaRsNS1w0
BfkFviQBct2w5kcbYaAYQI7yC68E5Tlk1JTCP/bHSFr6CaEcy3Es7d6nLNKayypPQcsnHhNerHPI
fZrKnJK/++UToQ3Bw9/w88TAd0oDhuLOKxsp25nBIWuAxU18c3v0omnHueWpOVXc0y+1FSv6hSV8
anwnF/lGSY+ff7dBK1EDeGOOSgpQ60YxcYhcsPnx+2uKfdpN8tEFXeixOyABsTyG153uspIWJ80O
cJA36YiDhjhAtjH6Xvv1Ggi8eIF032jRio66iubQXEI6+1d2w9aNYbFQurvyAJVX8Yyw6YRt2Ma1
z/W+eP/gBDSbOZXx5VHH8DKYA60kAm3ZVPGEQoQq1z8tX+yP/uX9geBCsNFUc/2pwdU8fKS3xUbj
HALw7ygAE1Xl33g/OhZUyJPUWsGePKiqmj4WPfrMUMH2aiWraZxpPxVJ4pColnMaGm8dnkk0QxUS
lhTOUpaZ9VU8eiBCJrVppPqTI7EFpS7n0YbPJNqFRW/YGBf4vqwjq4pbaUJqTH/DDBXwUJr0luqu
+AqIQh8ZQHeYGr9UzWB0A/JyhfZAekJv+jCyPvS5LBr1FddiawsmxcoLwND5u9asFOoZ7VElSN5Y
g55iD8yob/NADT/HBBDZ35ChR/h3xtfzIAcI6FOebhmfpaHb203ncPJzmloyGCF/MC0ELq+zrReK
v5GYNZApi6ZlpDZbct5M87x6+75PR0chcg5SIZvdNMBZ2V8535f2f9TYZL/ua00wPEPzPAei4ZAy
8X0hbokjsfRC6mB1+e/MCz2bDKvLAWQuKRWI0yDQw7xBTK945jGGdKfQVZzGd2mflyg6c2Szeaye
21uJ7tYenca7E4XHftuBzzPgwQFV1KyRPo7xdNPHUfj78C4SrV0nsXJ1DIZrcnqAHi/cSKocbM9V
w+IUBQlb4QnMN+L4q9wB01hHhA8YS2SYwp29x4RrlgOBmQW2Le+88FURmNk9puq9pOUTJsdwhhra
AGivsCWQpum6BkaklscZvdneWwKLASET2WXgYbE1k16JX4dc8D3B72vHRIg8mIoK7e89YAJpkPgA
HL38cDwNfrQ1egMf3H3CNwd3I4qCqbS9D/9yG9jTlTGOQ7378zE6mL216CrSOtVVEuYBPsLqkn5e
Q1HLXittsqUSIqnGOjYEHRhOpl5OPJyySmEACZCBbdcDVwob8klhE2nJ60yskS4oEllDkUeX3TWS
CF0WMrgi+OUlU0ScZ4nqwcGZWUto9h/Ob4/EPY4lpnCxU5BMAYnXA4IXCqNmf1qFIJ3o0VM9dgzC
sRQInQiNnKmJBTOTFzJkSj2RwoxpVz88o39sFXHO2ZbEGm3VqJamJHIf6P0+ASlWQaUaUv5lWrmV
uVdq1UhQS5wxde3V2NEOdBSsppYMd+EssNc4u4YK1WVMY+0pll7ObJBuXiBLxhwwt1kUoVSuVNKg
EpcQ7bgMomRVzZ2oKxcGf8YK5+gJaQm6qIYskIFo4T54y5P6CQrRPOqP3daXB0jdB4m6HK0GOVRg
Dz/TLmqhtb/2riAd/Kear6LgeCGVqcpMYpkNdiyrdNebrxwHb44z7ZzDMpiKeb1Q8Ddtj2kwGOlC
rzFHuzk4YIpbEXTg8aSz0LFG7mODFF+O3tpy3y5Cbbt4H3aOjFna043qsImx+tlkkD1IodisGZMh
qjoSEsHCEIUS0O210w3lRhrSFr2+nFyXSLLwQ8PzvyAFfi5qgn+4QaIOQ/0tHKZ8XC7CAQ+a23Rp
SECP5OqHS7aut5LfmcCys1K9BnURlKnOaOd05uatkV89nK1C0XmjdXF/0pTg/cJc1CS47vDmVEvl
hcVijmQGYnaK4Bt3ufnb2O0FSXKq8ELDo06sRIjYDofsLbfRS3BlHik11V5lSY8yLrdsl220ohtR
fJhgOa+SSFeW7QGQWellCuVlnks4wRIqxUtDZYPrHZd87QzqDrTktZ+hCcjQvyBXRKyaq+ZViJpF
rhPpNWxAAx9HOubsPB9YzkwyJxRtm1dIbYiDwvbKYtYw0FGACrl3kcb2bfOvqIjjYikLBdrTsepd
ESYLCxJmdJwEFWd7LdnNKQsWrx2HQVnTd8acED6k4zCB5tDVxGlLylC/4G3B18qvGSQlkpFJHKQ2
uEwl1f3w31qg1CXpETMEbMFKeUEvrlh/cYR2hrr1VPQ8gmk2BzzlyL9qECozcUZamgqh/J8zyOl8
ekTX7k1CtFfIevf+FPTDQUQIqtEl4D1H0jrDWts0UTJQIBCtKxdG3bSjHnYtcWOnjMYURpuNE1gt
0aIKwpe1cpezqXyEMqTmBiin+hPD3N4mYI1t6cyGbMieGQMYd2oLodBclMyhAoc2CON/Kc2bZfY5
8ATOlMZblG4N/np5rZVqZbObVe6Wd770T24aICzsOMw41TQ44eDNl/HYLZM2vuuU0pBiDwX5aGQZ
77dchKZ5owyuVPvcMsH03pU9Kq3uA/igd+27n0f0pWqY+cIQk4IK4PQHWwhA/gEXP8Kh+WXUU9t9
3yyUjU3mxbDG95T6vZS+m8t8gNXzxCGUHXpgt9zzCePO81aATJZCi8SSvphmvWYs4K64+MH+vycj
b5+lkYV2HrZD/8L+nRP+6jfSPCIsEXAwUF9+d9LUK1Uuk3iN0+MiIRmAtsAr8jOKU+C6axilNuqp
RNbYtLXPTDNxBrTKW8rSTTDGunVn7MU210KJNsfaFmuhlnokWIlyh9JPxbcT8GfeMF5MdoVGEXNm
s4vzyYK6kSbYn6qCa9A9eTS2Brc57Y7gmVKmaUbKo4HjlJf53JP4uaWeHopx9Xd+AQFrWBl4Y/p2
YhRIeSj2y97x3R+IZ6yKJaoCk0vkOQ8j/Mt0dwybFvDPEjlC1wM100n1j4Cm44aFvkmkOThKyiiS
igp5cYL7Eir7rJj+7E25BIhdqn3AfwywiPf3QMvv2yyffWJjlTeB+aKyNZ8RGRwnM0vJvqSjTmSv
HNuxHtg8KmxYP9v2MGKVVYAE+2NHJKapkxNZJQzJSYmAioumUVLzTnu/5S6Q8fur+umzV9lbXNXG
GQ1OVxwit8qJII1m3RYUIbRJ15RvmJBX2CiZxKaSJ7lpD5ZQ2BF9twEQrnsYYIATinSTnuPscgm9
z+4xSCa6qiYDXXoc2K9dOgAZiRqwatJDxjxZm54LxQ5visaxYNObW98PoTIjRqaHE1IVAGa4w2yk
0UB76IO00oAQB4wioIAJ5JfQSFxXm26Ww+1ThCqWbVyTF70CmDWOToTt2OJnwZH3TlF87yD5Mmu8
yUHUZGnUwJPTO0PsqLc7GwkouDKePBdx88VHL0H79lz3pNLSJVMlci+KfN8UhX8dbaQ+NZ0MEtQ/
lvWkEge3I+M0fX7bHD08HmIyLy2Qepmw9vHcx7ZH9k5Gbxq9iFfGJv3AZm1lHGRSQgI8eTOEnTqZ
BEnr87HTXTx97eQ2EwbenxhMXpcG5pedQsjNKZS71Zj6SqP+3nh0WarwqVNf8U26ZNIAvgXGPnSs
Szr5Aw75tw1EAZl7wMAtQ92YKfYSendQXm5kTcJEtSQveItYNusZl0p6qAuq6+idRPW00mBHpWa9
aWwbwmUWooYREzJuGyQNTssnD/3+djob1nT3XKZG+vNwGqvo5N2+2vckQgHavlMGZPGVUpFpXfTI
D4enCCjYZRLLMdnOMbfSZT7RCLj4ieLBh5zN3yAH1k2pIamcBHgSgUlR8YENH+yYVc+WSPtQ/4Zi
QCMi2AsrGELOmYKuBa9AfS34PiSTqxaFRHvLpc/wdkGVzDACJX3g7iD3h612g9eYbklRU7ozt+/U
B6/APQhXBuR5MSwGcVCH0hV8G6ZmbvGEcdxh1v3DOqx1x5J8RvP5BpjMhPUtb/ElODUQKhUNH6mj
Sfo0UAdL70+T20+rMl8XWcgtmkLjH05At7qBwkwzjs4tEbTx1oDk5Mg+u3RjDLwfisU/VfnyQTNq
pSCM54IZCIIJPWyf8o6IjJYI7Nivl+fB9LtP2K1hQug1eCxpyw5cnEsoPM1GA/ynkgg+xznhmeB1
1tWqCkI/MEHjMRLhZkuqK0kCjgTtR4B/8sSl61o4T7XswlYKeZCpRMoWivMzHQ3VGDtQPcNeQH22
UlvSfheT9F+5CbdJUR3XwNPw1hT/NxIDKWT0VVtIMabqPaOHHpxb32RBtm83G3RgLxzVGNKmDu1D
8RV36CbWkDg1zZk6GuBDtAdGlEsBcSjS2FnwMCI+NCxc2kR62Y8yUAoMXL2eEuJKhn1Hc/9wKo8W
FGdbkGKMNbHF3XijQd+uRH8QTeN7GCD9NLaj7jmGoTT5YMEqg3K8TiFq2aD1cvtu/xnF9zenDaAY
uwppps+fZ0LREOXO130H5tHpCeOpQ//5XWJIc4n/Rt+Yjo7nI3ZOmqi2KZ+BlZEbSkkYnKo6Raes
GpJMVLIayM2Brl+VS2rFzzfqXs0zsAAQJdeVvBohvrzX0E8goABwOmGG/ub5lTUHoQBCwn1X+dV6
wWJfE+xcbpnjyGx4wehArgYMjOxO2nlCf6JYq0LpLjCP8r/SonmOjUV4q7/Q1DzNENsnajasK6FS
gAqmaG+X+dc7PMI+M7780oNfxBn9Y+T6JAo3YtOpDVph2LztPU8TDL3eGZ6z5jDF+eJqOqyvDdpi
FV+JcGD5SV4EtLabSntIO8ZoqCVx1hv3f9wubj8sTyY4Qn3rZzRqp4dHa1mpWAKwM9pmDyxGfHxd
MKBT5CQB7B4OrXVnFTQRiVterzoK4Qld5FZh9U+QYuyRTp8IfSPzRS2zCC3rZIpi75Ki+FSqdy4I
8BxSwSPZEGK85j9h9jZzHsNhvNCAfpdDIebcszuw9KqhWf6KG085TssnrVUITstOfJ3mFE+nmuKq
6Pg31E9cGpEut/aL9Os77TFQgN577hLPGP3tkepv3TiDeI9BmNNj60GlNc4BJxmwYeNKY5vTScG2
VZEThN9lyzo+LXetxaR7CDLwVUpbClI2UxvVB8B6nZWKFTeX6bn0jU0WjpwWyYX6lkthlsK1d0sf
Wh/7VtUwXU1f5XctRS7S8LPSR4PS+86Sl33MlLcN4Lg7ng5CtiVwLKWo5kK3OlZxDJXWwTQZWUAA
wzVQcukrttg9WsY2LOIJbOcvTJIIvAq3/v6hNxtKZcnQI9T5Muvo34j4X2VR0DKS77qOXMrCm2MS
poTTCFCBH6US+VHBvn57uWfOMBxbY0QXIhs3q/gMuJwkz/5M/c9FJ6zUZVxJu/8Gz4tnDUCyT17L
z/Pd8mE+s0o+33Y6zpR/g4ZLFeEFTnXXl9SQLgOIoqodjK8wTYXzWJXur64JAeGVB3y9qzOxwqhX
GrIt9f0SqtGBUr9fTE9yNzp+f4tJA5yQvzxX1TlkXxH2K6gtr1/XqmW7anm+yts4htQ8mL6OaSxe
jXwHzjxrpToumIyJPU9rUkzJgWvKrmPr3mQ7SSsn+fxyIwHb40eQNvh3jaa+5r7+I+2A9A0qm5Gf
SfzpCShtzpPG2JX//jSJUiH/ffALTtkVGvyX3gi0R40ykHgjoa6ZSRjn3/1j6FV83TeusJ6C8K29
lYrp/WjWOamSaDfgbTrbUrx/cAondYqq0AxT/2nZ9oMG5iA5A/Haj1g0T25rCMGHO6uunL3jGbpy
lsV8Ww8Ao7SzA8cp4BvAgHPEBJ4rTIdx5Fpi6k3ZlD+O+e40nTjwYJYPIMqoy/SwE+Q0RjpJJSXz
KT9YKc1x9deP/akRaHxRy1duvopTGncxunA3TuCz5MoyEw8bm83QL1tF+O1u8A/C7K3ZZ5US7/O0
gkmdj7Y1tT+y8hkElYO48g3Lj2ksQ1kiF0LNXhJoqXkFDB/sV5CVY3hbDSid6NJSCZMzIcduUk2w
wIOnL6FAnpNAc6x8OvQYPL6uKL7wEBGHEucHu3RXRxYj6VwWEconu0m15ouEqqRQOUK4sXfZ5Pf6
ZUinnX1mVhiNcfHrcfwig4H4vTo59KPSRHIDFcxPDe+mL3iNCM5soqKYdwU4CrJJdxYn4KpQbl4U
jto0Yq6Ug51xL1GyI/uSsRU3LOsI5Dl7fam1c44CBSayU697JttbhMb0Lx2UNC3t92u6lnfYIbAL
zfsGUeWnlCsuxIVqoSsWAwOJteUYycHQAWQ5SrSAep/gLF01ethXrOvDFHoGpQust2+SK7b+R4IJ
guspd/e04lCMm2PeIWaYo16c/6UzEnZ6pRfW2u6CS6Teru9KYYHWHFeYslWUBprWWIkrZSPfWZ8S
DXfBa2UHWh+J5QjlPeRlF5n/1gj8Zd/qbGNn2HU6N5lt3eoJZ5OXUcxrSy2SzeyLWuzMYEWZMfAh
D/os1GosI/Vb3UEOxQZYyHdWEmEzKckYqb27/0Jv9QQuS7k3FA6Szzw0lG6ogzJECalXNyK+vskB
qPKz1cvmZ8qs1+WAC+3i67nBDodKIImxcA3qMDnXC4sbt1CxHRt+HpMu6si2NnlffMLorMPuVo1U
0L/uurfQcZ5uhnhilMILjSJN84/1MMzFMaQ9EyAvpzbHlMM20BQSepjHLbcRqNVk5kRniSVlfaeO
gBbcW3nZSoFXdYlvlv8DQ/vlxO/u3gAZevXa0IvdBlTvSpnKomanX/dUT/0qqoMaKJUEj4QTenEx
DdOkCs1owpMS4CiPqUrycJamtecglGeL2atrokq5NKB94eTveaL7xhQGzUzSZNmG+dIZv1vpsjTw
bjXMBs6HsM9tef1Lre6UxhXu806l8dqNd4CMPKvKJKt4XkbxCjpN+zLZCff5VDjINICRmHS7pwdk
qN2zd9CB3bRKAb/paUpNvBKNsbuxpDLeFxMgMJvZe2TfLzQDPa9o7RNZoNhz3Y2vWK0TuhqZgiwo
SSH5PtWEPmyvP+EHgvePeRQK7Xs7lhnnmDfT9o79Ysdl5zyZXZhf0FXGkM7AO8JkFs9EtSixSD7E
CRkJdSf7LRj/sHoyD2bCW5JPel6g5y/wcYmoxbDp+ArUWDArnNklpWwKr8lBpw+iSmCkCAtMX/To
fTMRO476yhGtBObISk7HwbDhn3aPL3PHTSo8GS/XWUrVVM+L3aOnAT9p8Dbm46UKPT6eqLu0Ewj5
R0WNUck84Pj601YGpu3hJ8nAZiKzBMxAEBpjclKKwdg9CqvbS9DaV8EMbqLQO9lRsbI641y/tZsK
9tm2rxZQhJF7SIEsf0Tg5YKCb8E3DoLBacYXDvVa0u6bXDo66i56ZrL7ggTicVKuUVncCFQT2ufO
mUN5Tpdl5vEUBpQViQklJd4PM0F+STXfAYSsMKq9q3fFtothvMpSHIHeWub/NvxhgW9QiBhFiPFD
LHKiOHpA5eOwIqGIprkL9DybKrJOviYAE9GyTrCcE/YeyDBhrXev6GcYKRBf7pDx5anKp9o20nOy
AVXUmNACpgq3rSKcxqTTPWmu3mr42AFmVgk6IVSnsRKbeMSNfhsEE0nZARPfQWheiIxWKzzJ66s7
EsT+Yk5CkhMnX8lJeWfFOuSnumtkfgtApoOtvg71YTbJQY7Zl81uZnjhSojVx7y6E+Ck2TdamcUM
RZiQ75qEKsVAXkb1W/gZ19PnEO1sWWislMzwvNKB5uc8z/thN2O/x/Tm0wrUEgq8rjihe0OjXt/2
6BJbQeKNagD23B4qJum3bjwBEtg7YQNXSU5yzNG8OYMvg5M0obiu3bO9ndAWOy0pTm9NVb9VddnZ
x+E/ckSlrZoOF1dljnPa3ZYkcQmC3fUGZ4g+daZ29vVQ/cvmyeAqNZ5EkeUm9X+GuKnbi8hFhBmQ
+JHkvWCDPJ7H/FzXqqovzEBtxL1ocxZX1/n3NxFbvJ4Dqc3ABLSh5d1Q+SbIkDVFnzlkH4Ui1FyG
2YnIsqlgwtw0S2lwAGemiTmZMUFm8YDmRO8F9LaL0CnN6dPrYglgO5K7hs0/biTFZ2EEMfc28vT8
B5qQX2ivr6RiX5CZcOs5JmWhF+r5Rx5MK6wAmC3AFtVLWnR8yqrU+g91bP8FEYVq8eupO2Kksf6M
2121caS+6GoYwZ/RSxM32+4uJiAYYEigNEeg6pTRIs/7Ckt6tT7einn1nnhNL1RSMKusDM3Uu4c1
qW7EWcnon6Q+q0B8PG3ptgjlvOHoyCjE2ebMdeORRMCd82tY6iuohGtyHRFmKS6wKUPUEvXvNeC7
M+FEhfATW/plsKR+93wEV34VaRhp/QSy3fos3HFxI2GWHvoQxVqSf52YAkCyxDOFrn3UaTiqe4oz
ZPhwanovS+ooZy/WZpBk1Mb5dL2hzs5qZHua5Q+JVTpPQWVbO60NxF2Tyi4qB60BaVtyeb27f0F5
s/nuTT7rcG7I79hnCZH1AF7R8TcRB6qzw10uK8Eo8ZcVmovFeTMvxbPYvE0PlJV79Z9I0THpIxR/
ciISdXWgADPH/5BMsqemQsuLv3SO12PuSDGf+O6O4gpKA5GwrUtSaaQHkFQJT1qLFDjMVHSTDeSm
hktice2Ss+HTfE/s1Yx2XFTxvCqaIsxDvvATprmB9oOrzP9lVWt+HrmptVw7kwRw6WN9OAVXy/7f
K3JLnwIGjpvXMDxx6rw+3FwStttDJq93GUl4bWUFlCxTRbSGccIrZDyWMPsiOowQcK2034QEIRzX
bo+OmGP7vBu+jOFNK8/79i8C9ZpauSe5XAk/lGObC1oPSPCQ0Rwz/tOLaIyCnutMInDvz3MID0W7
u/LPjcy3SJI90b3ID+hXDuYp2/24MU6JXygS6g+/4f7fZSqv8M82qFSWFe33wpqRMoIO2ffNiSRO
gnwoLmhusscK6RnDhgkCeVQszsIInQ9Qgi064N+7xudMeiAhZKQ+WHI/Y5auvn/eLx7CdP4nypIz
GYOMPtJ5ntng/G0Ec/C+CLpPQe4+yGncl9fDZnOYLNcUO7JN0FaHTtWocko9VnQNbLmciMdgaTAj
9UAce0TR/t7TlVXlHD05yTPxHoLfflYYeP3FhQ15i4e9y7KzBEHUcBVRktEaiFG22klpsX8wQf3/
rBKYYJeM70OPbsMazD151MBM1qauEQEXqx2dwk2uDhK9mMMOsPs0hqkKU7mLOoZOTq0Tubg+EznC
iPGIsZdLS2q1PzSkBP/6gCyPRM9REcEmCVW9fC8iT47GAudSoPLj60+ZA141fvZ2FgPQERA5UbNO
GkxQmYfftPyRFAF5P0smFsmh6gw2D4HOxzfGN6N3/Xox/i1+jsPweIhwjMS7t3sWZ2hLJZ0B3AX1
ZD2c3xi3L4dhYKYTQmRbs4rlGKKUKxSATzDMTpDNnsAs1YvJdexUaJ4VaUSUKeX6oZUDqInD2A+j
8Or3uwZCCcAJXMw5PZPY6Zs+9g/dEoNjHpd4j/f6Poi/8IHAa2Pr+WKk7vThe2juGnHZwKQ3UfQW
fn74lo4PwfgAnqheHWbGOCL3ZO/4wpTrtfDs/xlrmf4s0quq/aY6O2Slw4Lbv6J2ZhQR0AMwmEix
TsYNd92xKuCnu7MXSDIjU4i+zljCEYcReFCGlVGOsT+WH2EHgiX6P9Y1oqB8bbioYy7rq6Zf8kmv
7BJzR/QJRIFg79eOZUXP6vIVuNHanhYgJuPQwn10fFkfoOUHiP53sJOy5Dl5cJ6hTKPuEuQE3dAE
HAsOrTbgvC0bgd96JDV0HkebZGHKw8eHbLRIJ92cw2AUPQh/N4aDN6cWMyvCt0tXeZtdWCeuA4fS
4tUgkIukR2t7Yey0chJyu5vyREIVnv5TwWjS30HD4QUfdLrSffMW25yZbrKg3k9mOJPbQ55Sq5yc
1xkItwi9iFOf2u+AU0oEi7IBWk7MyDGoyq1sUpeC6LqcfkerC24XJTOrBEM2tZs4CnjcZIMwzBQ+
1MbCNWcF8pn5G+S2iQYEv1OdcwWMQddxUHK6dBQTzW61bOnC8QAtONO8guakmStB/8z/lika9okj
6kndaMvlVk8FL4Pj+Sz+xpTDEUlhNzTwvgiNnuY5USmo+Oc5/06cNRD3xEz7K2MDREylHRuTQomy
7tngK/dYZXg1yPBhH2csue7W6lOXe/ZL77TAT5SnGkxPbUi7lINVMMxQXuKhDRgZ4q0bDx0Hxywn
xDcmEvm9wkRWLS/B/se0ySQnTqviDkBsgGKM3SmRizwVh4kv2OyCehzn2gg/cij4lMi1/MvTc5PS
NLr41zGW9EvlgbV49nh59hIusTI+u6Bp4QLSOTE+dt2qRUmGf7jYAUZQu5PJ3/bGEnyu3Q3gD0su
/j2iA41sP/0g8RzwRS9dKF/K2/6JwAaCfKDZaU7HP8lBBQwBze4uPeM6TZ7vM9Jy8qieAyHLpLSX
gp/TBgqQqwPOlJnmr/CDSW71FPAvBI95PX+FZeseRB642vBhFumWUi3bv+kHwaSIPTxRUVhOKhW1
PmT62SNVYt5GRd2oSsqLKQJxy99C74RdJJu72uippHhKG+2GBDW6YLZTzD7Ls1hVVuSfyIwmpxtC
CDm3X81gVMG+dKFSITVyV/FVJPjH2DD0y8zmKhzueUMRf+ogqWZN2fatEwoLrkDFP7VshbBat1iW
qXB8LHeNEjWVr0KW1RUZvqFXsFXz1yT/PwlOkqpKXjN0m40XK3fxLxvWt5BllwDdc9HhJUT2nGb3
U3bTp6MMH6tTzyOZOOHJTU8UJD44sUsln5bpciEvSb1xSwa4OSen1CtmNeh5VEXtknByS/4f2cgS
/B9KgkElCuR0fCJaHBVdPCWq0ePuLdDCWGRamFWco7eDb0ZDCgxkXS6D+C6mECBfb7RALK6zLQVo
HCm68w6mUrcN8F9lORzfEotx4yB6Ho9O5zblo1Sk51p1qhyS5O5yEYF1eP/svkmtwtsTfGF33swL
I4fg+HINZgJ0Az1jHgf2/OwEuLl/A2A4cLx7Q4w8pVzq+64mqD5WI68c6VFwMG1sYLMtmEra4t1s
wzIt41SrSvRfCM3ebaUyeP/rUtpCdtQQeCM/5+y66X9FYsm2gq9pXaZ1VQ/AKR/ggxeamrmqdVJk
FZ7vhrjXas4kUtDmwwBwm7VFHLEKi6lQWj+nQrdUzWmwXMMqs6FOVLZHUgNJ9zD+kI9hg0HAT72E
/sEuAW8X4422YwyNeQ7ArDe8j++Naih4M62laChahNbNlAJlDa0U3xLuBnFo9bmSTANKIpXqf1ex
jaOYfbs6I4tMvJD/xSOzuaLaSoIuaUPdMmjr1qp6RRK4GymnF+kPHA5QacfQP3R6bzEQIipqqLBC
AZx1fFbkgJIxcgF+0bACiUVYnFt9H1KW0YjkSHctyThM/U/4kwfjhb6Q3rvVqeEPNeLHR1hlIwEd
H1xqvFG8We3qDCvetr4IZiZaA9ykzSUE6LWw6/9PID9awLHYo0LqR+FshnEnIobNXrmZ40WDSC/F
MfuEvdOAdaHsVMnZh5gJ/4+y+IVU86wgMtjFeaPfADKIR82VE5yeuWpGoxYVlumtATPnaTOGOAtR
Ss3osD3ZAXrg245USIa7RmTMVsRY30Br09G3ug7zqXu6CiV1BP6B3CwwiW9kit+FTCdfQlUiSCc/
AmOTvNgCF5naqtYzLC3bZbeWwaYPKV/mL7vJSPdTVxOiKVZgmu2Tjf4DEm7SsxRW+WRl5h6yIwlG
pU5uOD4/h3OL+54yqjOLsxWzN1BshyAEzuN6Sg9zayY+8aL3EV2Aupf5hfM4UpDC/GHRyelbm2oa
DXzOp96/+3kpE6FBPs4fMdFC0WLCT48TUgoXEVQaEMa090aPomNLwCDscSodCoilAoHUYQ5Whq0a
C8k9FTflajR0qe7tqIhszq3Gy+XgP60DB+ZOYGKPSMo7pl+6FTQiH9aRSEIrtm4OR/0Pv7uEwD9L
fDhAN67iVq/e66dULKUpPLKMUAqmrspvSA+jIUHq2S7akkYBX+LPyqA5nKmQ/WTPMVzqLMADrxgk
3/6Yya7Z6h6HxNPv9tPIMC6wb6UKZdEqNFuFCJB061xKnMtxe74Gtf9N4dMZEePt7zSZpTd4t4CH
X/46P6GZtGZN6E7VN1laIOJwGEihhffzJjw7X1rQLHajizXE1hVGBQX3M34ViIcov2FQa3HOnAfM
cghWrQ4UM9RwbOPwPKn5WMmblrRYaAS2teR2sOKNHDHQIUXNv8NQnE0G0br+JM+fUbN7GkKHGd5K
R1+8WgsZnGNoX2NVKG6+3D/EbtqwZV7flk1ghwD8v3NyRA6yLnKm/9BHGFXMXTvML44DrKSro4V4
zPEuUSo6E8upBlZ/uUU9hEWlB/biNww7T5CU1jPdodM4eQEp0MJi8gzHvw57QObJSYG6k1qV0znu
zUvhm7szrrBdMHX3PB2MqCiBRfhlPuU3KgQUp+/bNmhq9DgW3ckFYAZQrCmoGV3h3lBDOT4aeSrg
mt4wQtEdN6imTI6VlPeox48PrCWL9ab0DXONDIrpETGwU2W/8W5lad8khpSZNsCFLKsjJZD6w/Ry
+39sJ2L1w3DT5fV3Ikiix+oJT47hfNyOSYHPedh83KmbeRCa96yhMXxuQpbzvdMbwKjtMqHZoHup
Px1KbaSxAg5o/rXK0UiBoxM4QKb3PfC+UzBoR+klb9rbV2lwbLWNhiHRdv2nl8wCs+z4r8kboN6u
Boa8iIrs3otzs1Ei2+dIKpnDGO8DkNToZuh9h/dhye5pAOPQ1jUec9mNeRkhefXk1irxAPVwIhl1
GnTnRarSbfPOq9QLZRUzbytcVL5HZ6gcA8TBoN11fUrupQ51ssUs5BZZxkewu/x/sOUtg8i47JfF
z0R9RYwwSeb2Ux/3j9I2zT5uRGMmaZUlkkJuK3kf0tTObe3EH6MHwi3nr9wksdMlmW6Zk3KGTv+I
iRnNTJVVdqdogQT9fhd6fYwQBm30XS7J3zITXYfxJ8ENHH4wwslHYnOzHq9slvQErAjWsyKC9SUf
jMQlkFlXdk4M4OZ97LX1AJ6+oYzCBuQE9/YCQkgL4Uc953RTwubMIFOQE82ep9oED9oW2R+HhC04
l94OXwYeoVIxojZF5OR+Tnbsx8tk5FH3ErmpthbNMRyy+RcG68gCBCAOy9fI5Fpkwp5HgOrmGSo0
zh0hQnxU63KiY8KZRz6GuYCqzt76KnYE/4+kpVi6YQ32nxKOxTEAymfI9+H98emQStNy5lQhrMjK
Bp4wVssrYmryijEWOZnQJc5NHaggTeYnmE4l0Dc+SikRHvIEJZqdp3L0R3Zv3PqD8Mf0+mjfWoN4
lAzRSD0Ttn2Rc3jpfWK7cPY8f5Q5ouzp1N+bgwqj9k6+r2h3d3TtQkHMAoHTR8KhEqlZAELz1gDy
MrfhEGYsCgB5N5TYcxtVGmhi6USC5n76ZQeTP0Jdut5en2v1Eod/v7J8GiJN9qgVqsv3w9tDEn8V
OSbltudRUJVnd9QJTigLDRPwrPX9jGg9j20ccwHKOQBBV021u+esKaiRS2pmJkwqkZcbaxJwLueg
yPLcaB6u5QMCFZFysrGTqEoKg3a7GoSG1BcK2QqHcgOYZUBX95KmrLOs+pILYePTBdDKLd3E+QqM
GJVckmOTv5wMozc+1jSm15qarF5YyTFxmIatuM3ZRPlDaSumsmrOCJKLD19ypDMNxXx111myxAKQ
M97KB+ZjeKCBpu01Rsy9eqnid9ktQUspSBBHjWJoVaRSSrJcrcANT8KaTQkm0KRlaydfndH7bTn5
mfVm/wfLjdzJcovDsxLny/1qVjRZvqr+LILGKvIm/dfZdicV1Q/Nkuod4YrPZ1daAk6H3gsYq6nf
PfE5Gt725FoqbkmTRoKXypOs+bc2gfirLgC+yH6WzFOw1/7FFYp5JWqSXGTI9IYiyEf2HQqj5kjE
c5Bl62dTskopUJU4FJ3D4iLhSrBN3BMyfA9yDlwuW+QMHAYpqTyVR4Qf601paq8njd4K9adEKGBh
GxbwHocgXZE9NvokXGgnYkgLLnznQtjK3+TaYg7eHnTEFs4q1nPo037dsz7H3m1DPek6dBztyyZ9
Vezt1ekyGetVILiz0QypcW9PHYT7AzMTiFDNA/eCZ2+/3NBjRjOmnROkT2QlO8q7g93rdt3mLZVJ
KTiUYm2fQzRcZNPpn7fVBT5aBXqEMJa5HhLNQf4nfKqdIylKPh0goBbYGsMwIlulsk8A5IamM8bS
0BXt6ELQsxIWPv7Htl7TFMalN7ZYNyEcEQN8D2OeOOrkLrEv1vIXcKtZ8iurzMk0JP90QMe4Hw1W
ugZdVRNFqa4Lcp9akf4ipOAiy5MDUSRCre0ifoFiwPr0YZqIdV59wPthgkf6LLkbHksXmsGjehSw
eqNfjMQP7sKojIv80gSgKuHv3FusMrQjfuLTafF+I/WKWYu9YS5SiyxAOQo/AKtiU7FOXbbKA2vT
1KbkkwfwnUFGjXyptxJiXUPGYu0N9cE46pL8mtG2O7jOhwX3l+Rb+XeG0mcDmpjcVXj6ohxcmb1h
Z5zE8k5tDIW/iY77y58Z321LHiy7qs5+B8Y3iUWHg6dtKyI49abEWC69Hh+QkniNUhEL/HEreEIb
vyZ81EZ6i7ctKp0Wxm28RGPyyDkAZqF6NpBQ087V8wBbnooqABaR+xoEsqUgk79Cod0Z1X1oKS6n
/CF+ZXPIjssKTTfg5vztQEaVWtvWpA0E5AWVDVzz9uJz5aQrKdG3htDAd39eN4yL6vGG3aELmRiQ
fE4r7QSvMmVlC4kZj3dlyZ7NqkiQ5z2kxwNwZQU7Z1xbz3yKvw43woXd3Iv4/v2YsZsNS9VIC3+v
IWg2pp8ILt7MceEAksh+/qoxb6j1aRKuWDHgjn3R63+xIiJ6xz7ulDDrQitAQRfPyHTuB/6/DyFX
OuuPvi3DOxTMVqdPcQg5Cb223Ir0WrdBQaM371vlUzzvwxk0JhdaYowc223oQjPss14EDK5ub0U4
+N6+c9MplUAeJSg9QgPR8wDUkHvS8aeHbb9qAmFWYZBJINQOd+Fk1zIAKAr1DFBt/mkNojAIu7+f
cPUXUwRr8gHHOaayvarFis4ZpJr8ytD76sQElsEnq9SaWwlYyRrWXyr1kFPvwagHNulWHmLZhcBd
3iFLw9powGXbR24vY2cZHDngWHqriBzTDX3kDyDShdRSsDPL6CXp2JjO4ynhooJnKNup0pPry/Ix
Ko1oTE4eukFKoRvMmWsjzH3BAwiS16CDONNiWjieuN54o/a7tETZzeEcKDALRser5+Tp/NTg6LsL
wMm2+Ku86z3iW9B8isEzTqyaO8NGyGo1ilo1UDnlaJ0OLhPwMHc1Zgkq52JH6az3nCI3EYLC7die
pg1GZDRmQFjzMphrDvF622QCE/wRjiQ31icnkGRyYJl45I8IYUhc6lH3Sn1kfDYSapsOkqR0EsNn
nOXvd5g5ppiqTxd5dgTkYCOGzlNvyj4qNidwAIOvu+Y5G9xAgwdOQHEskLoBYld6yMr5lEjg+2E0
bai+ll498Qcm5+p4vhbv89XO/E4xTo3Leh4MmV/ISct/yeeuj2yBbhRzAXr3K4k6CUShVb/VKFtV
05E8yZDJCCtBzrXNaTjUdCJOEiqZ1cyeWKVNC4NDO1jdbdksGGOKwt8ovZ9PaO2G4WPq4WOY3//f
4uPESapalxk2czyzdjcN3OXEuOZJM8G370d3QLNBERIGGxMCOd+vbfRiNlgl2RhXN7aLetDrsTJp
8qIotPfyrtIAkIfKPyh/nO37Yiw2UnC/lIG6E31HpDa0dpiYtWQgy+0vHwWjUn2cG2L26N2NSeFa
Hickb1AeNeolfabuznwQNThUZxLgt2djaXnB38gdwv4CPfNgjUFzP0rKjtR6I+zlqIhprO3uxPqv
ki/NwVKIi9pCM+OaUQkQFgZztV6xg7Jqt8fWNItTXI/ZcuPwtF5rTzYrzLWDM3wjW2KLM7+8h5JA
b6CE3wRegSI/5/8ps6tFx2VytiTGENsbqtqRdvwY5UpngIyzmhRlpSdsAKxSdS++MAHq9QlkAEK4
gOPF6zEV4Y+h7Vh23r44VZYCLVuqQMSLABz3v77yw7Vca6YKfS61o9a9ZvGhE92YM4oAb9Nbu+pG
Ou92EnX7rMjCiq0sILXuZRm95cjl7ZyIBCyYiYaGL8msMiAPoolwxrX4Yl3G4tIdE88AeEKvlpcF
g8CiwK1HDqe+6f5Rs8Pktbox1ES45aamQmEVRBG27Pql1SZb7EudAytjsK2lcJVwhkvzbP3TcVDq
QS1XzDvwhC1zTrDQ/nokujN6nY039C52c04HYWf7cXlvZkBCbTmUjlUpW39std4fApGyZAcbQ7jD
/rQaZvnFFDpJaH45IDMrAXVWdTSlO9ENKuARH87E1rqixaR9Kfwp8UrGu2P0hwpRa6CD105lP0FX
7dUKa+Qyb4CJyWJyhqLvpyZOZGIHL5IXJa0H7xMYekzavE983NISNY5EtRgwe4JfhlPva8wSj5Kr
umOlNJEykFGnxg6+EONNX2EhqK6b/DNu5b6ZCVSLeo8sZmKz/0ZcCErzo63l+XHe6BJJGa5yfVkB
qFENmV+yeiwxZnrn0cIpjpTAMSgrn9S1WKNYerW84BYFonrpijp2U4pu/N1BMj/pzu5WIbw2K7Hw
PV2BE7WF09DUnyJ3Pk/Qa6piMXWKjGzNwHPsFLsWKP+XhD8SAF/P1QuYoNh20XCovRaT3VydajhJ
lAMDmexOs174N+0OQYBpXp/PbCgmeKf3TpbuCVhPz6qhwYCGYc+agAreWpPyyl8uW147bq7jrF14
hLDLIOd8trDLXAstSS98aVlWoKIvnrRNM9H3YV3xXORnYfDv2B3WVLSJRHqc97Cy9S/vSM1wDD4y
rwUXntHRRN6Mn20Mnut7AOn2jOx7OYLRhn6iS2wqtHv/7f3Djcc9Ejhy1JMbTElptEwbYT+pZS5o
6PmegXssXjrnQEujn28noFf9L5fOAu0JbPUYGtwejrzcpX+vYSfaZB27umTTn1fAZkoYRAHhbgEo
wNK/GyJPTKjRx4GmZSN+hGij7lSEDpemvauW0vc4YU0nw6xZssGhjBWAzfSvucDdLR5iqvMLkafC
2xlNl5oBaJ3acCp3EoAtcI5ERY+mQhvGF6SQk/UcI3p76oB0hbRe4kKAV1uPF/bymEYpkfJ5XCio
CHhftTI/CkN7ypnl0WBkWYaCnIiTc94U4W3NqVDIKkSps5M1mCtzUeAxNYF3ERJCnq/03AdyPoM/
N9t7ZMNvmp+6E3mAkpC3Cr+aiRfdZtGxkLYTmk18x42e1fY9oNpAbgd/4gmU4k0D9VU6dKK2HeKh
X6Wc0NiyBBbXW0GvQbRe4FYVPsMvAQits40P52PGZdW5nVjxkdc/zyxSlCGo9vDkY2k5DZydI/LL
mg4UEKVfTJ6mVy3cl+jN//zx1u43K5RWEHVxB5O23iqOKNf2tR6sSDn7BuiwxcaXtmWmDh9PcmWW
PjkcNAnt73n96Zg0PjtCXsAA1GyyE56coYJouFK9lJj6BKEwQ3Td3O+I0d72BO62R5c7a0EpI4JL
ch4V8N0gVNPn3+vGrn2L3yNvUDFFTCo50xv7tczBCmpa6Go4Xh8mzU0Yb2JptgsHJ/Gi2xhIf+VR
b1yK84w+Y8ZRSvUlE4Xby6/qeVkHJpE18WzY6MCXyZ1cMzaqQF135aQkKvOjg2+C+PF6L11O4rj7
/yr67LQyNLeOJqZkU+B1F1f8kgIgXl0Suy4szVWhkoas43+IOKSelTc2zj9rYOAzRg01maF63mr9
3Ha82XkM5KyGU5ZgpV7m9JOMYUb6FpRed6cV6jsne7+gxwjgzEjx+XFWYF/PAi5kflIQHvYdEuZW
kDB2tZHyZJm/Ch7c282mEs+zMtdbnipFCriCi1j4MiwzDr2XFUZPwoQ8yc6U2SP/anTikl00Rgsg
iZe15YtGuDPOVcNaahoZL07ZgWCHWgDPxEmg/NBNnD+OHHfsXyh1oLRS4Qcyke92Lea67IWtBCW/
XedLB58I5TewGl+LpnMB4QldWH0RzMSVDmY0NBL0j8JXi4XP54sXQkZY40v0Yq0msMVN4hJ0616j
PFBAYKt3k42GGLjIcpbpCk/937P2meAdAwm4RlBXgUECmKnAfaS5Xg3ekUpOh30xMsqPSv0jFllK
bsIEPIL2PZfch8uLBRxxkCIDnMohMaA09uoh+wqvfRRvyuH39T/teiEmGa+NUVHuLgBLBc10DmwY
lfNXskoA9YgMat6qBeN+xvJU8wLrLBRfNOXaNo9x9n7SbpQbeRQsf0M9eE2DzMBFWkpabxiFJ50r
R6/NYcmFm10Hb8siSyxrdBa3FKaTTxunAbr6VBTTSRBtRqHNPmofi59Fdhpf5l110+2LjRgpDomr
vzckl1YTqM0OzlC6o84UU0Ovm8ioyX32h3hUL5uLUxbbDH7pYEnl7YwWOQCe7MVBDJFMNUIR7IGy
h/+mE+Aco2gNxIV+AO0NV/FPDdDNLzmVMvfueihQGYtZfqgZ+qXvuWhZNmbD6Udc7azBwnj8MUM/
KfOgYEG48r9BNyemvTPtiwWqwVwq/5YP2U+Vywd8MAlILj86ZdRHnKW/EfMMfLUAdxP3GhuhWx29
nUsW/QfbPZ2re0Jih8t3GZffz2/K33heXbOWRZpK+lv3WSawTdD6sAB/67NEeBiQlI2O0c89gINs
kYXYrfJYNvNsDCBnCQxqpMw+jssvaegO9OXZMJ9Y2uVyp7TwzqjxUsqVKtIkHRsPlmpYFLEgiaZ/
LJ5tTQcb8AaTW//Uk4lZcV0HToTjAP61D1+kfZWsN2AFNHT5D5bs7XJt1edkphiBJY3NZfttaq/Z
XICqjOleY28Jjm8bBS/bjrxIfO1Xz1iuy78qCW1feW/bUzdxnMeNwRz1cJ8+uYesOqO1vn7b+jX8
lmEEkNv49EVCPM41ZzPBKrCufxZte4lZDUdBAQ8zD/EFp4MIK3Akj/Ei+acOBHgZYDmS1oSFgnuR
m+BOOUmzmwNSyq8HFhBJ8gMlTMFxcZvwaHqjp7q/S8BMNGH8sctqbdsz6RehGLAGCfryObocHZUa
iYpKbUqNZS2cYcyv//ZX5OvbBypai8w4Lj8ew+t7sdWY78GNDfr6Ov1DRcgCl2h3LBEpnUS475Rc
5+fWAGex5waeXkioYVUm3KxAxZVahK8i2gGA2oS+a9fsbIJb2z8c1cltWIATnyhElHXm3vk1pn4M
5Ssr1gA6V7bhF1IdNKLyoTACrvihFz7BG4zwS2YIxOyFKK2Hzq5uQVlnKhbR9pv8lAH9dkhIktUM
ZTbNG2DNyL8OJINnHCyJW39mRupUkNTfpd2ZfZUlURoxZYIBJcp7A3jGk0vqh9WWVSkHfTY/tKFn
SF149tcDpVN3QVEi7xUnaDShJ+nPMBf4Z6rzn0gRVG98OUN0Y3vqNvG2gUlG4wK2m8N2HD4nPoIX
eoWzYM67rJOpuXTgU3VPPbKwMsricrZL4MRWYHTy6ihyRz1vizZlutYlfPdsk1TQmfm33r24uDq6
4P3LFFDU7k4e/o7qH+7y/6SwzN1fVmSJkTBMr9I4qEhb+5FP9uSdpOHtxKpwn/owshFLmVekyG6R
mkIGkmn8upHp5yWdN8+FFQrrx92kCcvO7yod2d0zpmeU4+r9WSY3JGnRceiHS7Ij6ZuoRY6LyJaZ
MubyQq1szjpGndMY6prQFVQOwm9ELvvUcO4RB2qIyTnHHkSEKNmYe47YFwCJ+EGt350hpewQ1y2E
W5Eif1Q6qo7vs4Ga9zoEjNXhCGpiWaQG8sMplY/noRvvxOFa11Zwst9AnyCKc39IaF+qTJVRo4OG
V3VsHrSZ/SYH8zcZk2uGB/7oUr7GOzbjWs+LgFIf++VWCSFjAmUjr5AvCas1jIk7lHikTrhH89EB
+YxvuzrisNKYcEJWI6iZq9NJs/USqCyfGrKEIWHuUNpvmIBtfyeWYDSXHut9/1LmccraGCA6xeIE
B3s+xrP8+zyvwHsjb0hqC2YpnnhwjtXoOMy7NvW6X/yghjlP58wvEZzAyll5nCgPTe1MzEADP2+P
/qGJJ7dN4rS2v/a4Cf2yKYI8qWHTheTHkSsksNOpmI0HwAxtR14g8GdxQiacTHi3DvqvVBNhjvUJ
rZcP/wLj6XnO6UZXdscyiXF2ail46Sr3usTPI/r5nX0nNNAQJIXvdFYw47YL2DJnabgw0N49WO59
bfMXtjILgY+SKfFSVWhurCOlbgJL+ncpnYnaVXMhv74LKr+KLWviP3+8iu4SQ0zBRVUmBLgzUKYc
py6MunUvjR7bei51/L26GlMK9fGjfX65xNLjpwGCuTmh7tBz9pqxRpF5khofjpmt6fcvMVxmGhI3
7QDFeskO1mu2bqT6e+A98hpILt3pyU2saljVswmYxOo202oAkZynDzi+S8o2JN73G7cOLVkCtWFT
irQP4jybGBZ9W0H6pS7bx3NGH1WhtKuweQ34QwkAu3tH+WIjRTOjKrBtSJF2ZOcEE8XaNWJwW3OP
PCl08Gq+b1qjuJEJGj1VbYX8rLRtQxdLnVQk58RIVfxIubPn9L3KTGimfhNtybdGwetzbn+cWAka
IgrVBtpqPAxza4HFLawdtAVo7iaJWu56mWXL8MHAj2ofB425V/TZkuVRkl11dlhbi3mKVvp2PMDW
zc1bnPAbrswVWwnzNuFe8rpbx69W7ZNVXCMVU0O4G27KKuwWVL0L9Ubrs9AhpNl3KpW2OTDjMtlI
pIh1erOTOE6IgbHGXGyuaFZ1bnwkeFHlSm69/zNZPFCjsY8fM8QlQ6M5pqrxYf50WwXneXZeTx/7
o+Ce5VQD+zXbr5QuWQYbZGb4/RkXLJYs74DLHGyfUxDZwft0K4FddClZ9pp62tuWZUlcfUWRjBES
XRfujHUQu75WvIYI6uZlKrQgbGxtYZXK6K9e6oaS2iILeBIGpj8FJO4GAOtZpUcazleqYk2o+DCS
WC0W6zb9xDvLhJcWrWZCynKYWYJLoCbN+BuL/gFfEqBP/K6sbLx2lJvtW5I/mt7JXt737xqY2L8o
bE71+ztDxChnCOwWu0o7T1qF2zRtf8LdjwPdl81OCJL1FleEPyR7PpMP7fgwAEVa8jTfcW/DuXfc
FWFjN9c9SzwIarMn5e24+dj/hQhhaVX+CRrmQ7XyHnwvvFLmjqk2AHDlY9SpExDsO5OBcw4mzBF9
eRb825Tn9e2pMHxLheseLSmlKW+FhiQ0jNDJXC0zA2FkI5ZmTai8vz9+WvT3j89RFOgUcXFzLY5N
D9/VGEzQ4bHEyDrgKokwoRvZMMXeOlvjaC/kH3rYL4Z/gdW4lKmjX8r+RxJc6TaAPIHOKpx83wLd
f1ij0YfLNmlWI8PpIi+cBxn1zrqNt+iSTgJepiCjvj40rDOFl9KhpDgAx5IxpmMlbg11J7rU7kzV
cCUpYv2hEFunTaK8TVDsLGYXjOqgE8nopgbzFRq0wQFzaLosjyhu7xL5rjUrqAdzAMcrvY7iqJUA
l9ced1CxwLrk4Ih9t18l3QNczo6gX3EaqLIqUXH0YxJfGndlZSj8NNbLypqYJP/tIGCqdPw5iwzW
fwYsTdmGK6i7gZGMK2IfssXHbouNq6/kosk0sVyYCmtb6PQ8AITQjBBd50a+AOaGkIiVnfpXkdYt
lLrK0E6VuXsJo04VAgH0RU3ijXnrd8K83vtn929rLCY1Mox54TuMpgES31Lu9/BxY7VyxLCyI54A
TCyM9BzVDrR6VjAWYKqDRqkbLZcvjcU5fENYCuHmi1VWNRBv0RQI29avoXcmzWvmlaHrjEqxe3qd
5O86p8HZLgM/AaFt4x4qFPxuFjhoH+uuYPQSP20lwY0UP65vyhx8T57RbLUMhrWSYH/zw7lcvIHw
kZVecaC5bnV/hLyc5+/uOjjLKK2lnq9KhuUsvayM984b6KEyRu9jM9QTBeDVkavLMe4bkB2Gb9p5
afsqyOYzkCM6lvIGOfc4Bnbsygd1OGb1TTNwsxjIKkA0sfRHiktJF342rZTRRsvXieKGNKIj2wTo
gWhRC9s/VcZkY1mKYI2RFSkJmgjzdOaLrG0rky6Sn+0ihOOb/78cd61gDcpiuFgfdccmUJKkjWxF
KomboyI7Q38h9SNphFuD7qzlIxtZk7yeMptpE4BbX2AHsyYFv3lxbTHfgF3lJZIyCHqCpWtyXNL+
NPNmT+2mtrvF/7GkFfF1c1BHlBekvi1TaV4D2d/gGRBx5XbNX3VS/Jjv5S6wp1u3dFYWUgsLvRza
u0eGOenIP818e9fgO6cMTLg92la7RglTIYBQEOpHdjE0wAVpY81ckT8BjCJYvoPfxtNsEPM7zBZ3
0/M7+cFQJiz6LoH+jF3Ptr363LezoOZu13hJ04/xr3y7HO2yzyH5Z4J52JGTxOkqVVdW5ldIcaCd
jqPzUjcHYVM3T3xy2mc1gcTKug0wH75/T6YbTfGxr6l+YUrzD0MFjYt4eb5ePtGqj3vmgSuzFQDU
Of55VSKPffELirD3jvl+Tm7IfEVjq2lLjQ5z0NqsP3zZk5r4XfrlkKDybI8xBp3yPEYIe4nQ13t9
+RdGjQl8Db56qCBOpH0m6ofxcyScamS5FBQErLQRI7fPsX/r81hinfgchUFID14S+NqFBeR7lERy
jnV0SjOmRDjlrstYJRnxS97NcD2MGItJfk0Cxna2lX9UIB+1Vkw2724ASsqA3asAe8ci5HgclTdf
nFUv4hTs1/NwjFoEYtsj8rDD2s49RlLLzSrJ7+l5yTsZrWuH1txWVwrhETDCFvNELUb7gVYVA4FX
KybZ/MnBYPahBLsT4hqOOpj5UhzRfU7W2RTl9MJL3E+cGYPNkuVShScZSXlzJY317PMj6gARSZL1
trlw/2W984iSQqJhPXWS6nDcPVflgtRhdD63PusVd7bkLQuoeKTST+RUjDeigGMqoQUWJ8inPvBO
VoWJNO9UzUw0H3+FTkzqee2rolrwCbvdGqZa39IimHSDiaiR2FbJJ16Rk7uwNysxo8vq8HSUwX19
FRtl1s5GgCUqHFEm1arJjY9y3jJG4NY/hT7NVY9isVvyOQ8Kblfk73CWyh8zwCoImY0vWE1Fju2L
4ta2RrYwOV8gi0vVrVwTCzcnrOOk5iRQbO5BSZc1nvfTPD35f+G6rRmVNbvXg0s7iWmkXkEoI0Gl
KKWMg412ZIqrH6jGw0OkY9D2YGES7tU/ibsWm82m3S2EAdWMMJ9wJLc/idQ2CNwkVctah9RXzJ+p
/l5Cp1GiDv77DY07IQA8+ziuo0qe7FfZmMqkgSzcYr0mQtOL0m+6FVEvH/2rmUWqeYPIpc3EeEdR
HyjWt5g6P9XCT73pv2dT+yAGbIwPnE/ywZ6mw+pwcomV6G3TLeU7pPv+R+SE+sWwI7fwY3NBLMIZ
LQ74v36Y18O3LY5bsUTCq4E3Xb1bkdJKMtZL+y563mFjl6Onmgpn9D6+dxcG38JgvbIj7rhGBsZC
N2QlEcRavKBBHN6kI0ZJVJ8hCCQs3zfDyojUUpcVV4X2XIkjNRo5y2G/sxqyxM8wHClE9I2FxJDs
/1O3eMFlEU8XlAPTIWQKesUR3mv+kqBv2YpU9BcB6UqcfhetoDxGm9zpO5WnBFn499WPFmX+vqh8
ThDlsQbBVX6nrCmIgC+r2yYXXMRkOk1/+HfaA1+zazo3B8XhRTWgE/k46VeurKkwh4XZzhSboV8i
74uB7hrsbbkzRi1GpwDRz7pDtseWL3wG+oveT5TkdeEQkWA+MNY+OzSHXs0v7hF3yw6xt8IfiuzV
CCefDy74U49oPUlbmPQWBph+P0if4Z3v03PeY3GC/J3gLPzal0xqE6RfVyG3p9Z2vwradEetwKhy
kYNLuZfmH1dhLMD6R2/Am3GGOIAZiJ5GZqphG7C1jrib+2Sku5RiFUgpaiSMGWu+0LLwGUkA1K5g
gADodL8IHkdHDivirtwt6boYmp9aujorVCEAnJH3rEGr5V3/LGJfjtOUauvELDUg7qKtB4E6VmA2
klffNwEWx6BZY8/oa+8FzrpmPhAC7m4UDSRemXjHnBPBixb7hNMI0A2TaQxpP9hXnzHgWmEfStNx
E0iLoCGWiI7BOvtRtAFRYHnAuRUZ1Swy7ynsiwAkuz3wC44zxDogwbYZsX/++J9xgHG39OpSJYBz
ZhRiyOIB7oPB1XWEZ6Q1H+EmaFiQQghL03oMVBbXyRRIQbXsaoWp5UwKnbwkDR6uR2fc1u/b++PM
g+Csgm9UAObplFlfOVq/GuFaILwjpjhDc7Olhhv6eTGOmzwk8v7xhXYk4VouhSKhCKMauRXcxyM2
LX5gBO5Y+7V5AHMDoewCEt/w2b0Lb/6uvW41M085UcZgI4KygwfRNFgZelXrEQp7FIPZGdZWYUdK
3g1D6Rnhk9RpsY+s/7anFDsD5TJQ77sD8B962H598dEKcACgsQPJz5eTneSU7pAWfSRzGqI4sKkE
NifWgapUSZlzT2FEeDGZ3GLmDPuSiayAt2eDXIVNS3/xfZ4w7AefA6AtgGjjMAMoAQGePaDyxv87
q3g/GbkeZpZJPs4ITKNWGbBIdz+wO+HtNDRKCklxKt2sxM35j6Q5ZNmw9vxqIPO4OvjYbt1gkO7H
bFf+lzQt3ooIsjOXTru8CjVXMawFOU2tDo/A9KnnHgAJDcGCMyGr1AgsC4K7ARu6uir9CzXDNdNa
sSyXcXKI/XKfn4nESG4TheXulSDa/Mivd81d5dcKW73mW0XWbIlXmO7Qs95BHqI6KC8PpIbWpeuZ
C6DobBzgFRJWIJq+bl877+INlqloECiTcu4+u/LreQilZGVtg38oQ9hHVcpXGoOJ4kETJ0WtbsF8
g6HfwUkDs85izbK6M81sG/am5ZVCXBsxC6FlDVSm79kFWef++fe+s5gUPDK60IL6pFPSgkWBuDWW
4FJQMXwqz8KYhOJsgF+UR2WDWyWlgsCcIOyOHwCnNTCUMRSh76CLlau4pUaQFBMpfRf4x0B7oCcJ
TtMFcpDnOB5xYsPPLop7SAHRDgC3CJPGz4WNxNlu5orN4la3h4CI8HOC24Zj2l5tXhk+lzMW7DM7
kXXLZ+2HFj6evfXwEJb1gIUxMYgAI9ZTSCapjhywSjrBihAtW+RhrClyX9dbhKJBsK+IhDMNqYm8
DfAAUCJFHsqfSpFLM04w3Zqo3hNvpd6qOILaKOSL0iq93SEJ+/K+MrGK3ti2WDN1PYteaL5Cdsid
0Q++QIVqQFmbvnbU1mQ6bI21Tr9KyuV26yY0ClXzS5l5PoXcvOVJz9D3te0DojVd7i2x3U1NNfie
G8rCBAXKgd/9mV1yWRz9IrXprvLzDxUAn/Uizp+bRhbd89+hxR7QWllQ7WWbgWEuf3XwUJnlyWK3
k96r86uxVKo7fzC44GHbx2pvIOKKKmRpOSABbONE6c9dZ+2e5DTfVcMC26FlSk14Ybc4syZusGdJ
8gmdneuGRmjQQXqj/rnHZa973Y2sheqtgGqPIY3NFhPSuCdq+zqp2g5IFo5RaZ4aMOqvRkUSt9w1
ZuW6dMI1yIwxPQJrBNJPdfXsOdbighwvIg8Tbv7GEr9IDpUD7PxkJkrhlUEqZt6yPoZxXcH57vcG
SsCzi8i1vehY8J8ars+DjDTzWWsukUN4KNI8+o7SX4JhV9NzHQ6i25fj0dgD/QLSn5cD90duIhV2
NxvTHI0GcG/wmw4Bbk4XkfM6nq0dLkVjK//CGGPXyNvVVRfVDdPcN1yePThUAD2CytyFZJRRXwp6
tzwMr/n+RKmphceNtgFa+M0lDWRq3H6Ar8rp5EYKHRJ6EEUpIBCHF4GLgXa/7+sYqLMybxfGHSqL
bn9HovlGlVa0Fi3cuoiHfLuWrK/Lxxj5823SEEfaQpGukDSNIx/mMytdXbehpmhBe1OOZl4FX896
/NvfrJyzBw1wnbKW5PAbD0rGBpbKNZBh4L9KbgdQmT2OjQKzKq8ssoMMgeg5iBruoW67OQera9+4
jGKXt2jVrYcflp4qdhHHjMU50Q8Rtd/8WilGfaHhH6azJvypJciC3Ec9NVxlbBjjSZ2IB0zo0pbY
ToyL2mWJL4Mo9xaWsFhXKW07lHLhxR27cOi5Wq52e+RtmXkrb1jbdNDImD9cEM0tS6Z+dut6ffgs
ZEPt6LqRZxmy6TIeWBa2pkDCxd0YgXOCCemHBkQUi065AIrQ2ZBHPdpg7/SxSTTt7fto+Xs9NNTq
LsIfU0EIy/zAofLITa+OPLVML3IemoKVDmeumoEr325393XCNKDtZhB7WHb1FfaH7oG2u0EkVA66
+H3f1NGxABc6S0qkEkmK0AX77sMeX1HWndhQZRgjlgmpQCX4xzJQ3jGMFvBuye4spMG5wxtjkExV
rk4hkM8D5in5PAyHX10KXGJHTSdMiRqUV9O/+jyFzce/ZXQHFzpjrqowwQk8klK+bi00G9mTVclO
sSxG1ElZw8NaHDUlS5t3vI1lUGYTFoIJFKyAEggVFc6VEK1sur64ZsJCbQWtF9hxfEaMjycJrAuP
92Bwa33gyXUnsBTmp1uvG3lLmg1Cbpmz7bwMjD6MD+1P5mF3KjF9KDSPrf/DwE2frLNfdizMb0Nn
C21VpKwZD0WMBGN6z+n3Ryng0lcA538NC8JcQ9Izdhk8QdSydHNRrT5bS21ZTnjV+xjt4WYmgMdr
n4HQTOmM4BWDQQGwV+j5eQ1Hy1EJ6isYKLePabixzd7YPtANUlEubIcT/HWKlQvK5M6TFx6dzc4W
RdJVNBDSV5geurE5W8K84zAzuqAmvA+GLEkIQVRcz/pEHsEEWigWMgHpEYXgYGy3OTZnuyuGYFWc
bdPtVwQIbF6gaxk38k273kP9xce9OwqvMfn0DjlIJ3Ing720ND7vXwm/6SBhhD+1blRSdl0YjXHT
qJUUBg2O0bu7l7nK70SHpevzF9STH7MbCKwPfayexJ+sHwszkzpYcRCSdbQrcCSdLxLXOQJimX00
JdZNEgU4CZ9GWtcvSkxp7np09JcAwq4NHjxpxA+gB4ZJlFNOryjoXK3az0QV/LY2Z8a0r7Nh8go/
vYMcqAFkGL5pc+zA0UTOGmVWGtgZ3vJn3qCUF6eOfuGNL80X6nFCY3QytiM9KZVldovO/Y3vY0B9
jF3UxZCkopvOIMtp9iJZEJawkSwuG2Isngs9ZLrrqvb7fAdGV3Cio89zzEIW+NvTk2gzNwFZeSkX
R2MmdEPi+zwtGzrA5/IcTa4jkhtR10wQAEW3T82wotZ0NEVyu4YGe4zKbYWxnNRvl0AAjaX1efUv
9nN/g1+S92w+Yr32Da0YPzWPnuRzw07PexeUdSPqa+kF5kGXeXNGnZma8b7uF1gNRCPJugfMcSLr
Ul4yTn9UOLUAUfWTD1m+jng5M1Rf1cOff5j7e9ejeokKtclECe2/6SClV861mDLgNZg+UkolSxug
qEBrZvI7WF/6ZL62p9qs2r0rIfKBNSaKrppb2+Xrcv4RKOioi1KpwrJqtELA5A6rZTpO75KLJQCK
hdOUerHBtNL8bv4LUVthnKfQZgG9/VhiQNKJfRl09Q55aAqWQRAEnmAXkk+5HIyflYS47Vpu5jD4
Uf9TfzYGuG1Frd10Wj17Z7tyiLXh/9AGTcDoWVpkyE7eG7PdCBb50QGS1hKn6Dj2bMq3xn96JR4j
BKFwr6Z3Ux9kHKK8hoFfGRSlQYwKNAhvNYxWwit87+eGeP6//QhTA3BBYUz0l3OriEIcjY1p1tAK
deE6gkSpCeV1CoMMF8UUPiEu7P0aOSHRHuKEyU8XdaDIx8a20OPdRGzGN0Tg2nrWCe/IB8ESCsCm
f78OiGuOwno9Lbg7P1tvCd5425GOC9PrdSLbCHkKCtAbGzODp7CqbUiDeDa0h+12f1iEICALBQ+q
YTsYNa3ODxBXmOOy5IONU38MOg8nfsgjOBvqLQwUZpSs3Y5CTfqNVLI0l7vcG15dgZogQ2mMOrea
BWAhEoxbifI/bfDcAbsYuviOkPUYb56xHNOs253Z+mE8Ll7B7DnaxufRDvRQXm90wyHis7zL5fIk
MFI+3ej+ElDw4gx8sj73UIPmO7iOnLSk3T5saZmPDBgQjaLtRbIyjpLO5G8xhMyHV936Tk8DgiM4
cEFVlOEAek0AagOMaB1bGnI9YlCbn2ZI34wfR7cp2WUsUarROyGCNHz+zY6ls36n2+4b/mbx5ojl
knH+wsBpPRqAuDPsEAbm5kagvjedu3csuCbmg76YGBPPBY/6WqPvKWr+2xdZUhv3Sz/D9rKYEMxs
DN9Y6TTQHOS2thGZWm+T1zCJt9ChLbK2R5o3hdtgcG/7XxbmidpZwYI+03yL2C6lvGgNX3vrufMy
MX9crXrcOiAj6TEwBW9oDNbuOkPfrYtvXLiNWQAd1RxT0j48qFVZau7AOXzJaxZzunrrzAkbKkHV
wmhBzu1qXnmlDCODMC1k/jrqCiGJiTn4Ij5El/rEr5O2g7KhpSj8T/0pBP1emB/3oZer1Ccr7LyA
AI7/E2GPiXn/r37AOLj1LsJFUQgPxQupfhtZ6VsczvlLJ8XrfdFvX9V7uWVH7SntWd/d1KXb9eGv
qPGDUnyRTNEe0AWOf9ml1BOTJFXqPnxlVnfVngs4SxqPsUaov0Ja40VqFyVaeP/sdypVFxiydXwX
mfjQSyz4RVofigVCDXgUNDqRfbQB6L/pD3qMn6+muVylN3qpFblp1JrDGPivRvM9M9eEoudDnaAG
1l2olmEOv/cFP/lyQzfsoCdJYCIcnToDZH9S5dMot4EyLsWBgRWZ4u9Ws6QRcwOZH0Xq77hSHDXS
c78cio2LqILkpxBV+1upn+prnVPxQf5mFj2hM1l4FiOOJVxmSqisDpVsmVw+sr69+bGXjmn3YuBJ
OZKBfxWz+Xo2NL6moIiT6uaeWQyQ8xZNEa+55aRg0duzkIry0UAFzXIATqTybm3sLDFYrnZ+aMBl
NRy6ZrvCH2Nduz1iR8qksqofnJIwbIrPL9fxd4Nr6FCJo6+021MfRDxTFrP4Qgr3iWnAzDKSpUMj
nExDoV+H9Jy8DG0PECelr/DpDyj6k3YQOYNZxKBEAWs5jHhaKmTvEWSKY47Gpip5FowqQjm4mkU+
BerY0NMUDm1+CK2RY5vr5sUxtv7eLCguv2ll/Z9cmXvUkSo7S0ojPgejwLLOYijTbHoKpFX8HZxQ
LZvBjXNy+wiDM2mWGtrlcf4mXeTYyW3lfmH68WNs0+d0tq2r1//KsakGHmChZJKLWIrzLh3vCx42
ubKRKb2ADi6xpWPX18/df5O3U001w28CVWjhJUjXZvO2jueXUWLAzGeDkrVmGA7jvYLg7Yg33706
TUQzf972+CmrR+8ZybGXKwyCXrK4mOHHHA2IA4mQeAPjC4gn7GLb4vX9p3ZKx5xIhDc4i5TX/8G+
mgmQnCkg66di+V68oyW6Lx/XcuumATc4yeA458uhv7P12u+XU0DbYuLYV7Ru6n8wEKmSDzVny1Sd
1nZPNJFKiYfmhLPNgUzWbyONY/b2TTa+gWNkmuHXmjhW4ETDPI/xodVh8FkEjZC9Nl3ulVNOTgFo
oizLkZRvDO82/LG/tvidOWwVIAT1Fgb+7t9/dczqe5LjsTkZWD3oLWfsFzujrDmXcMAi6U0MN9gN
JgAYuc3JdzzCDvbxcZIQB5OVRlfGS79ex+0vj5znbOMNPqdOiaCWIv8O8KEBUb/8xT+avSEOIEsl
DQ3h+rDDJXfLy1JNz3lX/eFp2em3hia5u7QqcFR8nA8A2gz236yzMy1zIqXM0hjhfk4fFGQKifVE
iD5YRWHnQtHIywZ0+a5GALz0gCbqfGO0/ZUX+XKnZq3j1F2yqIX5y9e/umR3bjXDlEa/pcESLVsx
UVZ3yzpNNE2uYZ8LPMr4LofFjV21bn6xCFMuRMY6ZwkCt3QNef8z8s6tBxhnngElVvME9oxVdlm/
OjoqyfGt9F6Mchp1tLurJmLlAqbnz0brp5+zPGnfATAz54BqEmjx6pZe1epnuGnW/CEpau0Nvy3y
p7MO7OtqKH6vYMIFLF+sV0RkFiDKGzjVTWTH88g87FfRS2SF7vu3YKO9k3X8hK52z0sHwXx091o/
6gHBxyTlXEMpJIiUN6Nta8zf8tSuu2qnAh29cit7hNtmnWTzywR7t7X9WMMNqHjbl2LXHrA6g1vG
CuGxQUO46wkSBRPbpMU5cBf9LbYHoxVctvl9ZCHSr4xmgluHhmHp8y6pAcgOHLqdYhgDDEQGOiaR
r8wQYL+yOJaAuRmS3l6e4VauANc9M+eHl8nwCuFaAZKFQDBFfzUJb39RBiUBYnMntxlP+/2ekVOO
LeKl5uQsmP8QtR/AzXAlHGhrN173ZQDaOeq+FXcUzjK4ePSOV6scUqssY3rtlzI2bN7aOuwiKh/3
t4YBybu+JJY8UTKFOOQNHMwQdIFX+gf6bG5TfwVOWybrYv20JRho6bFjCVPPoksCY2Je5ygeDGdU
/L3eQxMAlYxJwV+fxaB03iOjebHWkVdAS6qmI7HqhgKvlMKeah6z/8zDqoXC0J470K7J7/M/tD4/
lh/TrePqYqRpx2BlWCMP0BukcDSucd0kii4yPfeXh2hWWgE16dvSpd2ej3mUo3OkAoMwQrJulphN
xuEcNWWGuE0RuhzaW3fxvJPdAFqxH1gJNcE/vmVLgoNWi/csGXINY18AfzWpO1WrJNnW2NaLwHjy
F2Oy37YgsIIU3LBLP4UuwJI4hRngigLTaK07PHfetXkQCoCGw5ViwZ17Ec17shKzo7+PeqxuysP/
gTxoO8iXZ2XELf/vel2gW21wudE2HXfr8wdCZXr5vaxsP5+NrSHCUtNA9jQYz42imIuRaejcHzKf
sVe70hGfLJgs29chCw5SHTgmG80DJPeWAXpt6i+KyyzY/5dDkiPitdHel895UQ076DgBIVbarz80
NRbaOCrg6BidEJzVOnaUGEiuh41/JiKptpQggozIgR6Hwb9nAKw2Gom/DM7h70umOIow7pa4VyfW
68mTn37I2fvyBU7vts/yeWLLhpr1mJQHHZo8FF/TUO8nfnJvcMZkANSlH6kKV1o18FpyFUayc51N
+msiOxEiLoslnVmXfI393irEjPhNf9ySXI2l1XGQiaaMYS5Wpj7CfaXCLgKVV0h2pUdkVQz4krGh
i5vrn3h+VuKdURH60Zs7Pf9CBeXDtg+i0asbDFrDA2/TMMdEYbGIpbXN1qYFMq7Y3ZimhhXPqNtx
+epgvQNbBNcUWHfSZLEegNb2NWV7ZgdSabn1tX0KUglcYiHoMWO470j5myxsyVXxZhWUWT6zaKtm
olrwLn5e8pXxFJaZ0T2pNEHiTkurFnyL0U1QqlUYdKRKmxKL3A8biKJvOyeHLh98fXZKOSglzNXF
QZwb1xUdWUlYojWgPN8ZaA0zIQu07WLSsE8NiOLaLXQ/UhfaWHPs1reY/gQCwA/yBWTSHupBMxte
dg8c6AdoWRMLq0P5J2OZ7UnK3eqyv3WLq9IUnwI1dDKQsgAho5zz3IiBRRMgBbEuXqxeQTip70Tz
jEZnDtRRpYD4j5q+/YMXkWpSZm6XLIBgajdM1MEc71FXSJUjvri4B/cEJ8n4GVXRXQovXcdDinSq
tPeJGkmKPt1YxNfD6XY4vjlgvr59IP64LE+kBKhF71ByWS40lf3f0b2kan/i7ZVCj/7V7h/z/zab
B5Za4qTqNMDNIthluCk9IpozBBEh/PjK0wajW33cjNrtUg7w51+AP24rltS+6nl0Wtx3LnIsKXD0
QQDGEz+FvL11rxDnGrYg2aKSsGrncY4zEiYjDKnadfq+i5PAEnoZz80/+fbwSsshaPiRI5FTHbQW
60CFrmSCdXPNOiJZCMxLTQaUhfOugDx6dxUDBjW7i+dQGUPUEmpkOwDjxFdydt9MCvK1TFuauZ6Q
wi1oT84w6J6A2CfXEmwN6BPm57qJxUzJ5TiGwiY0AyJzji8Uv2W7fb+wU6HnFrx8mUiVqwHNU+jO
BG/GSSRVkFBEoMpYrCCCDctgrocnv6SBbpw3myxvRDg4jGngDAe4MDmY1PGy44AjJIQELE8ZB1O4
eeIZeotBH6ATqeSUOwiva+E5Th/wggj4iRSlqr1/aQ+XSqXf9fqfQY5w4rq+ESXC0tettQfVBoJw
uN2nmvul7N7FcPxAwHTHXPkbDcL3xsgZLRo2WXON5WkTPbMV/Rc/ENIBLrRoMIJ2fnkjvJYZGJeM
HGt0hEWg6D8PBMH2u0EA1VujtEUxbnWysc7gFUhTGPy4yR0d02P8cpT/v7pSlcmCGGIVDyz1zZh5
UA9eOhbEuKrrIlwmY00UzJtMf3d+GvJr2KABNdE4yRSiH/rTEM/2baj4XK5ZzM2EfCufBKTURBil
Jce3WWArYZXIVZ8lrWG3Vuc1rC2mxVvhxME9UDg22faRSYJyGgttQtUvxdaqndFhIbwdmxC5xHCk
LXa8QuTstQ0k8cxiEOvFM6jXnYD1uv/6ASCcySNjcOGIjECYNlOfkij/gbmM5TDaKmk457nIrHa6
rLcva0hBex0ZPZn6jHVgXS94xlY+BOxwoKUBdklpTuuHi7isBcex6bjrQr7JyK2mi5XQeUixPvTx
isSHg12u1lUMHSZkCulMLteOB9joHd3tIyT5mTblkdh7X+Ssht1MMwkRsw3DofLyxq1HUYM13HQj
CxxIm34d9+RKiBD+Bj0nqxuMrVufTvkgx/zHF+uK9WiU6p2L8APTZInl1veGob+hZEwXVf1oTW8L
yNSxmD/EamlZyRyjtEtg+kXzqGib8bbgIHCfUhVwpGvMX/GtwbTsE0b6dzlgfDsaaGQ0Ma9SOhQu
LxOSJzv4v7r0+JjjkQ8Zsub9/Gb8ZyLqFiju5I/APgRo4AmxfvHXBk4JcWIKB3+GCfXaAiXiKTBX
TSNSPsvKlgXILDy6L647CfWfEHwV7p1DQYjl9aIlmAOjNL5AuPwE2Xy+dVR53Gc7ge224Fc2pYpb
fTA9+QUgQiUdHo9Tk0ZRd12I3+uW5hh21VhSpKmw02o4b8epjSMkbQ837tpLtwcnwFGT20q7ox+u
LftVoRKlIhu3s6e78NS5dQUVG1nYb/my5rrBkaGEFAyNpv88YRlf3yJtAi5U2bxcvgeLuGrUIxtQ
o/M4yD4/iaTuaonyiPfIRihWrzC4D1oLriyLvPNsaH58/py9PAmS2Z+X9fNfRvNBdLqlt8pLSBwr
ZIF59Cws4CgO0n45jOLkcgniQwnsETScrqcXWx1pKLOnPIqR4V4ghbwzKyU1eHREN0mR2bUyC5L/
TfDbP+1sHOGctC7/rNffkbOLQCAZXCUKf5b8EOme4eQ3nrSKQY6QzbZYTd0tMDnEzqst/Ej7XbqJ
MiyGnuuo8Qa6vlvJ4C5Qo/vzCk7E8KObdVBbdJAGXPXOLapEQc9zCT+I172yEHzN/+ml4H4ulMEv
qy1YuYqpjTzyxJqXYx4V1ZjsIQr19Z2dUvTKdRrpUTUa76S75ZwQp1cQFqsn7wd2xekh1r+qyMsq
I2GQ/+7M8OCURtq+gBQPC7F2m36eAU4yBgiKlGiA3xbkblLEyI7abRr19vZHTW0N+ee53uzTnBq2
9uZ7G4q0ypONVBg3u1DxZ+3JBbN2zbWJrOFM9+KyJxVoNrQnBzGKljw2doo0KYBPLSsx3qasA5WD
VI1uoLLe07UTe76lCA8jr7i2BMRnfGcZTGlBQWm0sq09QwuqtKPnObUwe6yjqtPcVGdmZfS2S42W
b8wXpU8hMwAv73L6X/3mszWGyNPChByknp0Zzww04F/KTLvb7h0vFOU6cgiZDLvivmr1C3o316F4
ULhv9IlEn1FWgDkD1QmvYkRzts/fi5fYTz0L0YuNNHGxoT+MmI5vljBKjXKckYsg6j8p0ayGFJHs
crEpkb+YoDp567zQDsxnPAH4rjOdmapiPVQSqQsO0DL5DGlDOtXsDsCZUm3Puugd9P5qY1PlFj8W
tkA1DecQvV8kMzWqarj3RUyI1IxJOj9xXAHwT/Olc9/AoTIqnaeBNFysETuXVQslnHjQv1Zzifr/
Qt9yq+smjQqXDz+Vhj/CwJL91mDcHh7Ps6aUT4Ui02BaRc8jOmF2hDeQA0ls0vQcMzYOT1DsAntj
II7vuDq9yYpMQAParcHwQjR3ljRSbxJEcm+FKmuWTpfxYnPp0l1TMCS9xZ1LeDerygFNq95bm11H
DT7hZGX779wmj3qPuoS6Jm3ReLaNfDaKwfTqk3JCrXeCZnJDGBoSK5XvXO0DevLPEXh2lq4l3qSH
qOWfhfhhsi20C0DqstxkJbB+UqrU763a67BNkBPdpN+EM30nNu4KAGLc5hWxdBWtxiPCNWm4TpOJ
os+4HIm/o3wpzUGcSa9DPVxWvCcJesBxEsVOrwgZ4vYQRlRiBxhJBdJd85taTaZwoAzi4VwlYMUp
Qdc4Rxmx0yoMA+GjkGiuH8rLjkm2Hffu+wAzdpLdY/Hv2onDz2Cn1KhxLlZdzYTD6bifk0dDjxqe
G69TyO2b19Rw3XZ8RrANAqYc+YiGL1efY4Mp7/yedxus9R6SX0jm01wQkbvr7j6ox/aXk7mM08C7
3iLM8fVyv76pKCCe4AnSl0awwqthqs2e52pM6ke3v8DPgZ0e81vSOT4N5Fp/A9uXKoF2axbuSzYH
igDnOCXE6/bI2+B0Hxq8oiiuWpdNnbcCY33et/i5h8f6oS4l+i/IagBp3ELpNThru9Iab/LBzXFN
24cgG+5KkusjymuQOD2QpmjSJOJRVuFU7mttMRPxCO6lYCYK7EE819omM7gonIKb1PtR+MLogame
doYnJcqTPPwE928q/CcgSc+zBv4qUHGe9j3t8UYYzF8q4aPFVVzRcVIkAFrtdK7JIV5jqzhoiVLN
myfjWDaxcHeZaIFhz4jXat2zjPtI9WFc0fSaZbkT3pZEdr9s12zZm9nRQ6UXYSeJdxL7arYT2ad2
G5OSoSwikA4oSDDFQ/r1EOpRkvr69QPCkXq8MODln+AzJxAdRblu4+MipRuDqOd5AiPVABtTzmfS
vxk8eJlf1mqAXdoPs6ubTgMSmrXdxLNPMpoy9N9hYmpF7rRu/nvmgzWcP/dsHeVRfFmk2Uz1rsi4
9FrflvIwtIYLkJs2ID8nhRgXssMXKoE0+77svbrF+aGmvPZ0hIjMbageecZ08rsuoDiTv/EKgqe3
ABwhJ9X7rZtDQg55fpExqV0F3SWQwyK/oE8lyhBC3AYLrotcrWmnsDS/wgj0KTqw97a7ptOQBTga
OTosCi212Ubfplhw4WLbsZczUszCAYYCV6tDCVXBdRhZaCaAi0aNrb9589zTVOTxV19XtRGVZkS/
xW2g1aMtB0vl+W4RUkNHguv/ZAOYSzu84Kx8ztfacuPqbMKjLKM/+5yaPZjXkj/2AI8IWuLDgf+8
4PqYoermUVtfuixU/ESpEsvf+HFodcZZ/W0OF5O6CrzpDjj0nie3DkSMHnEEjk+PF9wKQwYVzCPD
2WRlOXSy7VViOAj+oQnXiPi2nC/F+AL9eLtFo6Or8ghjfQuBLsSRyHbvHYfQjuUw1wrcqEK3jY5g
6oWMasjwFeIZUn+qAjmWNe4FJzz+mJM8h/3gvgiCOxD2XJ1Y4Rnfyv6e4Fc1yXwqwDxD5tGe/pMG
QPaAZnA+rRhF98ho1GzckiWWh+t1Mm5Bu4TWgwUd7QeC6MiAqWoNTlZ3q8+w1R4o3Tu2YhUDTI7s
chofHLaVCctESoqPkduIJKzQqZ1ZIkIhYUmG+c9V4jLzDkLNmEa4lSIoxvVg8672Jz3oH+3nX7Hk
c2yzEtfeY/UUA9Y75ailcTLrp1+b+zeMAAUo6mNoNqoR8JTSX59WX1tEtaOMdXnDMSzx2sHL3hC5
TZLXlqayy8TjC4cZfGFJ8AzRO6yUd0/QGdQphQPGQavICQJ7qqDRnsmooQuSQprppw7wUiXBLMsD
vGIfGg6u6iK3UzOOveKVXc9BMVM/L1DH4Ng/r7XWvLpjGSbjWUBRRGmUuRIskq/MMdg+I9FFzR2R
R02Cl/d4DYxPRBZHqVVhMAZCUle29B6lAsNn01LT4cPy1X41kMvo3Rbwzk5CLFnaA/nTgATpFAaJ
Zq0n7ih7hWBhaUnXEYwI6FIpl3U/aamsUZ9mitiQ35ShC4boT1Uz6wp8eQ/8PfvaTve2lj3jQDt7
05orrKU+cfIa2dJqQXytHuOxEqDZ2nunxROU/daxSQpsrcxa86s6G0CLobX9sACeXQmlcfGaPRDh
TuhMIba1s1GewMbNbqbHFMU22yDzSGGrb9GyStnSRJDsWPp0e0hCkKdxPFl1ggQscmXff1jEsjMm
987T5KZZZOubM0rE+FuxzWToobiXdC0uW84iGDPoPurxVZ6HxvjQWvy8Pz8V4FZmlbqXlj/zTgqR
A/FdIqv95NdjVzJIEVuHkkgG0K9bdkK33yBukevxbYlYS1459PKUDWWKFEfO+QMyiggUw0iztFu2
DrAnorJxFWgvjiv6oA3vr+OK254k5rPgNP4ioUTwqwxyCgX2WJu0LIb8RviLqOEMADUqXVShpjPm
CcOARb1qvTZ6sC6lNaqjAz3G4wEghM/WLbJfz3qIYq0U79kg8skLEEc+0X6TV3R+UyxC6BbhT/FF
B5UMcTm+cW2rW5X9I5BVWmZNsMaa0cgD4vrIMDZakBVkJ/rSE5ESNrY0MLIfZPDwsoWCBtebqryj
HCJ8/nuF8BWSB/GdDnGrt8cM7YeL0Y5bhNnpxZEZGGWiz9cINjeS0QABwOqZgWoVRE/QZxzvOEB9
vi3hk4ZKgMsRq37p/Af89TMfjWnnnA1aT569JjDpnBY+iOm/K9h/VhuYQYTyIZrd+yoRVtFgwTKz
v8w9HtbevCgm3xSEYp3cX1a6hy9PUIGnXaT3cPLJ5J7ZRitUOoDU2OKpgiB7TtpaukCkx3GtEYHn
c4SAy1jckSde7trSC44nDu1bLfDGKUVP/B4/kjtgSsOC1+PSnb5VtAhRIAl0S/+oPiYgfiCSxo4D
bSUX4xUiDlU1TxE10Y5XRGWn51rI/z0p3LkE/yXuLmkejy/75IDnqe7TpYaKLQuGi1SY2BPTElsx
lDL+PWrGzxBeAbGlo1lgfG7FeF2gr8Z6J/qqRLQmqXE113VhSeUVNKxb+0ZKROOG5BynmoQTM0mn
CQnU5FYYKxgJSUq1gjLz+HVWLhLASbSDm3GoWS2wPN1/sggy7pqQ6D5Jlfo9fPtAmHPGf6RHUkpp
TWZDGzqrMFekA6H4fEC0FGhV2PFVIYA/kNutxU2A432bn8ioG8gn+o5oaLlnk7zTfLaQ/qKlLpCs
hIcnCjfp1v47vwvK2Hp4xNEWf2pPJer8KFAd+cGkTK3WZWS1/58ue37SoMkY4kqoANFWehev8qg6
KaLc1Wdxpg27ggtuYckQfbXsk95FGtMKiZ5FZnBmZDHyTIvm2BlhzNDY+9H6D2DPL2TEKNbYAAUL
FfzdN98oGfp3JLXtRYAOnwU3xJdygiBUOaK5ErL4OfDzGlLvth/aVv7/PBdFf+VMR8YLdDO0ehhM
qD3QjbaT3m+TUgUpuv6X6tEtreKIt7MiQziCEgXQ8Pap28qxCgzYc//o2+t9EHDox60acm7+7tzY
aQ63UE3BdfLHmumy50dK5b8JC2ONaJMhGaufLZ1kxm5LyHz0g6w9w51vIN53QCzyTrS5dzHgghJy
AD958cg5SO31C1PmcYYyoVA97xAuMQ6PcZ3jWxSjZSTR/YOALPPpFngASkcCFYxIR3IZILraSZQm
WxdBLSdQ1F5urUYvVKzzEHFcsdFkHc5wguVZjioH9CxoX7UrUHny1/4EpF5uWPuJ2YsoHVn70TB/
WAA+Vx2wp54ypMvoikXtD8eAiUJYbdD1bUX4l5ixXw2Jh0myXFRx58XvZr4VukBfNnq4LH2F0NkY
c7uW2iDFfb1iofFEf29lKlXTIpEJCva+epmkDqlRJXSQJ38J9qauc5wI3Wj4briU+toy9OD0hDjh
GE2Y+pBjKVeApw2vuUvT++agHk4vIZnN+1O/z5bNxSROSdJt5IH1b2K8E9EYNNrkDU4V5scOKb2A
XrTKvO1RkCXRbyNs3lYSHtUHFjxu2oP3Wtf9kOk+pN3Q9pYS7J3/nAkPn+hQiO3SRnP5KqyoFb8o
LVdTrT65YQ7pgp3TXCqxc9vT3iaxa5msDh2uWJ9GrO1vhbP4AMnhUb9UHFNHPCzOpbfPrTBy8L/4
AkjqO5LjewtluaIqwvozvjxLuM4/QSzoJ5MPW6h6bCuKH2WEVPyu1dpn+2+YJggzaTeUSNusN9uQ
7Ebzr0VWGXuk+t6NrzVdwNFptDKadFn1ud4PeyEvHZ5xa4AgvS3WPwzcHJ292uVe6lLhxHcbgUI/
dxbuASfCQW3jjiQn70I0TjD8gQxFTQtXFbDaRT3er1t1oFRqVH52YZf8APhMLYMDaPEaU8pzyeXK
2K8feXxT7DU+UiB+aA7+0PD1hw7WQWa1JUP8M66IbXNEg9Uk9/NaVrlQhosceEKLT8I/YbovZ4YG
yBKrFyZr4atTxs1LytxbwLurkGtnBoLwjCuU/UaGeRyN8cViki6TqHmeP2kJy3UYWRtDoBGBAgAz
aYdemXcgdHU9t0b0Oh8lV/q+QsOr/az0xTYeVnU8TtZ4AtsHHQIUnRjU2Mh9AaC4DDMPcpShzHxw
OSZBBUhEQDnppGOAAlnskB0SkAebixH2zt0Wk4moNn4oJ2cAE+24FkK0EHrO39y75Y0G77k9xzOO
9dibdVqchgAq+zCBb+77kXpbLIi9R4/4DCxGsnnSEfAR2tk95yz9IM83020xxYSQoHHHyoyw5Udv
gE4qDRwj5AqduPXQhjP/sNBzLv8CT+C8rfWmq32YQ1nDTp3+o8jbpEBsUQ20TMMB6ok5PYqVWjOE
ikzbEnsqXRWdMxmrBKRJXOJOrBTb7/d/y6yQ0QIB+kT59KDFemIFa7D1q1naQnTdFco0bzOFAJmz
uqphrKXpCAGJTHLUM1PJPH5IjJSE9wUNdEdwsuaWpbFogw7qcqJP+k2olqekyL9bBVDTOeOyZuZk
YY5W5A2V2vbpg9wxzWcX/BnkHLVsehgKWaRAjiEILomf3OS7gc86ZNuNO4bWT+nyX1gxg3HMhnjN
TsGYgnslq/w4upJntZmHnCfI8aXsXARdHljEzp+6fs6OnlnRgyQHgZqj5UyBCTIZnUgSCpTn0x6u
CHj/ZSQuyHjCZiXhM987onf9vklRpDfhsW0Us6bbAgY/J5RawsaHMiqwzZg3orynNbZjWQnLL5CW
VfBUlKdvQNdLs2vCbRlyB2J36/jZjvhW4KPZVWAQjjWBWHBZcnfkyxipK+OZQYm02/neJyos1/X3
Y14aLO1taOM09lpKsU6CwKV4tmcdZxgAU6yz/vPEwSlELwbnTFmR/vxil32iec3Y6vk1DCQvWTVn
NTRRTfv+0ce0Da0Plin0H+9jObcj4au52B3TkE+aBPMcPkmXgeOS7Tp3DiCtQrsYXebGYpKv5alM
Ukxp+BbIKQTAFOHqsfaNVS+o1LF9J6Kbd2aOGNq6aTK7eIinsy/DZOVPHId3Dx4kFYsOHarrBhBa
D25zE0uEU+s9yaA6Du6S/SoaAYcw4RvErsrPcPk/4KNphMIjUfYbTuW5Awn9E+zNXMRgtgHyKoVb
GKDL/As71A4U7r9XswzPTWetaBuMmSnabtR4YQ0BquMkVLmMf4CjjLUAPv/mqDX9I0oyHGM5Af4F
CWr98Leav3zd8e5nCQ9OcDYANiQL2zKt6JSjH6XqS4IUgtBnlL5/HPjOqhHwQxxeOu4l9dQ95DS/
0dQwUteTO5/uvtPBddjF/6KnG6OzoWUVKHrBUeUbrIwAbO8K9qjmXLTld624dIa6EwNaV3S54N7I
kZBxpjk1WOl9mIm9j5SYF/GvWLwP2ODVE/YyseKZ7ggGn6XGtcm5IDbmw+Q6HIiNDF8Nocm2MxXJ
5B43ZXBeJo6BZBB5bAUUnE+NwLUAuQFB6YLQUN+7pBUMzWJwDcCR+36jMy21wOtBZKL2B+SaKOFH
yT2p1aXkgg38BEh0wbPt6bm1XupIrhQUA9c3u7pRXyITbB2Z4r1LXmXdv91QjFRenoJL7olgJHb+
yvycWqivFikJPYTyAwNCQKdg/9Ed5qh8VdQbwV9X0My9aPJyrXHYQVBslSActG6yPMeLiDcmT83o
0tn1PMztBnEdrRsPxS0hy1jxCi3h25AmOsp/I5bQRCjFilWbigueHj2Ar19OuFLxIULTEG4AmJXu
mdxgFG9zz7+FKaa4iaQ/rGRWB1PZljppHJbOhqY8TMgekyWmy39SEZBzk557QfqlTTLii3dBYUO6
WwzXPeSRpjtcS8Ks9sRRe1DWUcDHPkcnPvWTW6Ngkn38xDW2HJ0eBv9ejs4KymDsyGffzF1tCJ7u
jDDEvYEcZIm/yTMVdUefO4BgXCQUeNoVYhOSV72jmeoYWRfN/jM6UJH2oSvrHPVvQavq6h/UNryo
joX8RgqM+9HtmSJVkwk1s4bicycVGEhVY6z4kHz0aCiZA23STrz6+hDVr8XGthxDeunhRKo8A1XB
CUdY8EqYL31msIigqJqFXA+oM1oht2evUfs8PFm4ZNpEU4rOxxGpytSswX0MXG7f8Co3t+dZkiR8
AGweObdIVzQd6tofXUxGfpPd6j7t/A3rwMAU6+zG5oYBg0f26FeHClkO3MYWd2KM+HvddUxw3lIG
5BlDlLQY2evuqMakYdCbaLx8frj9n5m4PslhfOYHPRiDkbe6IpTNcRqJYTCNomQdFsfh9NEm/Ve0
ivxgehVUEpr3whjPMrBV8LtOX9sLejWsMASeuJWe6LRbdSRS7NlZ3tk0JFkmgfTUSssiUvMabiP1
ezG+0n3xX+XGzybUGxj6BRZ16jX7pP6dzfq6e3Li0dRLZGaVstjb0O6aX5hnkV1uQWNpS5aP76A3
iuW8vH60IwBTvBplQNYfzmYWlHlJVHNDT9dv3CE2igxJT3DP4H9UA4DycOwYVojvLBqD5hKHERPS
aflgqIWtQXUrr+YBQZmOkkGAwFsiRlIZDgoQlWYmdA+p8KvLvGvOgWralMTUSEz0g6heSGTyKsZp
FqlERVD3QoRn6gBuGmuL0fn23YCeknI3eEzbc6VEDCEHbfZkEx5RcR4WGcpNtyiPd0srxj3b4TCY
woJND7nz3uhfqpKpHiiKKSQBfAD7cBBtp7X3pq2dd7FrpKeMsJ242T1qNrF/R048vC2pmtNPOlFw
zTbfGPVRdmbF1itCgZ1L/9y3PbSNO2+ecwB75qxecc6REAyB9owDKBpkxjhkEm3Lju+FX1C5zUvD
wwVzc4JqRSuGpHNk6Z+rhhPVzCjwlgTy2QKzUyPl9S3GiSEqJEZTgdwhVMk766rNK5rf4k9XI9mO
z+5HFryiCYZ4yfqzpXjEX7ypXOJ8Kk8Em4ICn7Vm3K0PR5Svne9YScs7i6HSt14zJh41a0yo5YcA
ZRBAStjB1Hur84VF8foHC32pjLsivxq5oAf6tRAt76eBKlvOUnDyg0cG1HfvgDGvrzlzveskxIOh
s9Gd1TfvPxgUeq00bskKf8mIcJsH+zBG464MBeclTjNN+WBlOxR09I9tZEicrToPdUqYLIVhVy16
Y0cH3LLFXFPrFaBg7HExrHgcfNNzXfjYJ2tweJg4Oefc3fFZDiIa8dDL0ZtuSU+Or6TBPXFbEmgO
fbbtnDvinvRIUaFww4IbSz4uQXKgBj4CAmkhYJeGe3alSsPdObu3hH+dealerCvXdrcuXA1WuHoD
LMyHmlRVkT785eOeahRS/xiJulDldqojKVVu5VX0Uzf7sAF0KiktT1e4G2vPQTGLEn49T618UZ1O
wf3RkWqn46rnrwOJIK0oFcqUl1DD23B0PrkMH6OeaXzfhaQC3G6QG+pHfUAk9wcQuqCt9miHga6o
N8+hG8A9SOGM5a6GRLHNjQDBhnUzfVvy+m0rHdbaKX4I/ISkWfiZ7xStRYwwbZ0i9tlWrQylxXWK
24uUfdUdzJQe+xOY6VGJ5ClMfj3dN9WNv24bN2DKPUq/0oz9ViwxU7fUFhs1GU/RT/kJjx5Yd2Eh
bKIDKq4uQB5s4hZwqpgzM1Qv+WrTxm/AETxWi7zpTFjAOFAMPH4B3UGiyabaMwKuHVVh3QpTLIk9
6yLWYgy++D8jaJzCO8BxhyII2jOdqin9Nr7T8F+NYJ5dDM/pekupgHP7YLoVFXAKhwn6EiysGg1E
QbcD9PHJVlC85dZEFmI74Cpf92P5ZEpS2pjo8hxOD//yiuiz9+M2L69Hzxkcn5gBEAOfXkO1gkgw
2m5XREGQ+m2FcTV3vTYFZeMYJ+qsfGf2wvd4Tc/W+47Rq7a8xpJEzlnqcLA5cknooIiSl8daL/TM
ovYz7FJeaxSTmzWYSRnrKnmvlsgEkJIHurLMgJFr2CB1DEAhp0eAqw0fVDaN3oUDM1jNv515a29M
vZ5+5giZRDVhauI8TNUCQspCLmn9laaBcSaFd6pchqLAI6XmgVIodgHnyBd/ilj2O1tZgKSCKf/C
wJYS2tRN0+AwdKHs6YW4w8J9mlIMt/u5lzfbU7Kif8fTmuaYeaU2UvYvsVI2xLewdApY1oiZDTZ0
51ttY01EeX2TC3Sh1CH9GRP26AquYf5t+sOSkjp1BY+tWX5bb4KuFE8ktaqN3JOQpqWneR65ZVDw
R+EapO83kUX4ztw8y6O6KLT8XfARNU3X5ffs/GVzC163UUQparZgN5OhsKzxQCuG7Opi0jNol3R8
Gt6B4YeJojHV/3qh8k9JawN/Nr3HyuCEU/8vyHM9Fhy2IaUOkXNaL0UmcFKG3TvNVhVSakUT3wIn
Yr5avm8DyN5VC+7l3vvfeVJYkhKcfUFAJ4g3i5WphXKIm30dbCp8XBv4lZ04OnzksUXUMJVwQdZc
z3khHeEvnuqvkRpGqtynk+Ljdu3wrIBHMXasXIsRtyCqbYMJf3ruRJ02bCaOPR2UBb/vIjpSIvXl
Wzv5F+QK2ekJV/lbZPxgMVzGzgiA46h/ICCMA+YpFFGFgvsgSiSTJFUk8nKcs67gef86mK7A6i5b
88zGHRxAtrFb+ZS19coc8W0+hRvFpt4lyB8KZiOA0mcouNJ7iCDGURan5UZB9wGYpt/eJNn8u+q+
47q4NhIHpdrRxtObsuAlgZd4wtUiifPSoxXFYJnS8xhcq1QeWXfd29M9FMMmnfuEQCb0HYLS4zRS
Lcv8b0SQrWvDF6MeNZYtbMlmIu+OGtJ/fXGLainKBPr6PfTe4tHVrblSatqvySRTsxlneBvYC0zo
lLCIGRpV+1zzGHER0GEBPQJ+rNTYfHJE9CTvvcyCwestRxLnGtH+oeH8I97PejgELJbsVnWGs8gD
v170zjH+4TmHk1JZoEaQBByNMYj2RX4hxDh0ujAzKwP/Sw7Oq3/2hX/qH0gwCUJsOLviE0iu14Ay
a5O/yHDo8LK3kWv55BVh7wGbQa1v+LjAMIqB13w6H/CNCBBgsriIK9kZaHvCmEfd9IyeHqQCT8lr
3WrNWoWtEoicGcwOk3O0uEgNIdqKN0M57ifSi8Do05R6tGaQjOVQmCaMMj1XWcgEmZ0V9HQZY7Et
x15hZUOycu6O5db1UKQMKV67/O6DZ3qNmm9NlJwhp+vaQNMVUMfodocBsE8MxROmmW7oIZhTd7Wj
s+pmaaj2FE7IiJ9IRpagr8z5UH4WdvN++xDpe2bZqKielEFjVPom8zfFkBJYBS4y9vFQ5qFKlu0p
B6EMgiNovbPQxvyH2QJAiFThBgOYx8JePjJT//I/B46X1kigOrrkicNlGYqgawdezN8TizIXSY7T
LvcG1mUzice778emFdaB4+YeAG5g6RKViWnnVF/L0xSAVxRpyBW+E8Q2+MS9iXiuLNyX0fVA5ugQ
vljPc+C0sYqAAHJ/mC6yQIFrN5HJfzm6MuR2BCFDDLfRYjylBFjjt90eNCmLPDfRGX9SVvM0mvbd
BmvcjzDpuiNlMMrDCofNRRANwpDUu4vhzrQKXV/3pH5dzvxOB+xYZa5FnfFOdWflnrM+PTr4DddD
NG6UuliELq3WPJQgW8ymJffcIxsIdoOoe38jVcEivnayQzzOds5327txpVw3UVOGOkidR7W3Is+I
cOwA0Q8w6HscOYraIySN1gDm5/fE/EFFvzbhYhX74m6sbZwYumemVaktuyGlrsqh9Bcm/+vT8ymb
TsdFB0s23RXLN1u21Owiy6A9XiG/FJVwt/CRtmRtlD05x0Dj2f9fASqUSr8vnnMHSkza0cyf6LsQ
MANq4ZTFD6Dyk9qRpBCMoimYlLEtENxxG6m5yje6xemPiM9E9f/OQ2ySx/UBLSaTyECWaAIPLGxm
2GnRLN2WIa8w1m3rchpPqbnRy4G49P7P598sQ2ywH03T3No/8Ov/vtENfYlZWke82UgpEMsVfVb3
g5ZFfRnAI+oYW/CHZ9/NAF7gv8hWUZAqnvBhpbkyCXUUnIaI3OBYFabNm5b/GYDC98lcS4SVkkGJ
A+SNSm/WZx7/YFtVmlfFOMFh0kSR0ECthEWMUjr4WasLqvVzKUTM/eQ2qB+yfIgV/NpX5n5x6/+8
EeBY8TY5kfXjbPyZKZIjxkWnJ1Z/hDIbZbQlhb7xassMeOb9HVl5//KSWfv1XY7H9OZdQro8GcBF
hsZrVptgnTww1bBmeAm7uwkmCPsNRkQbVjZeKdYyabHf8O6Jg8Zgzml+ylpzy75EB4vOesKvy4Fm
C6UvY4PoWOjTqpDNXfLUDPeEidx/OeKBbMMveu6PWa6LQPBlkUfjyysv8NrDr7vCrNLJf/E4l0kB
Bro8qNiciSxbiiPeQ/OtIBEE2O2A1MhflhycaHS/vF58FzgS7sAGCo5a9e1eH7eFK8X/n6zTf1Ay
ybCa1FoDAVETNkfEr5QCt9VaRwlz+NPCOuhNpBAsFVJUG60GbROjaZIQRLLNBR6g/73t3CrOx0le
C9zoIDYv0noH9KoU1uHPatEgu/Do6bSxbDsN3VmkqXJxMcgEqYR1j7qjJX03HSuKWzAfU3K9yz5r
Ez5Gy0jEPru5lS5QYvYE2KPX2KknJoGceLRBbDWWotU9snLKnIGOmBbLFo7UlB/ursPZ7ZIKpGHT
H7LWRzt0P7cQ7BIN1sqPnZ9V1VgehVyrfC2fzjzjvYKPkSJWAZkNjVCfyauBNtVJaS25Dfq2SYHa
hBijOG0KcOQ25X+YLHIRe2NedQEx78I+29b1+OE/Gd2Ek/2nb49y+Us8qv7b+Lq8KVBjCqHpuwTJ
f1li+x5sXkgdgB+252KYF+PpEk7W24OiKjB5zaxN+PbJzZZfAAW3sgwU7qF0NalLFoiQ0fuF39Bf
phZTEebH64wv8NyidOujzPrxQG/nHovzQRP5VzWMd7F2HNlmyI37slPC4UfhiFZCRyj4WFlXqoJF
JDrqG1xSNw/WrQDY912sO9FyzydT/7SlJMQMZQfRgILyUbe7Q6l8c3biC/oV+edx+fnWI2aVUZu+
AQxBk0yB6y17tgpXL8OGvcgDq2Y3BfODXvhegCW8JZJxDMixCcexg6n/RuY89TuknsUAD1rGCupZ
V9/g6mk27NejbbILgKtjN6Gm5LEvFG+CKg8RYSBOGoUf9xk6IJXe5jlGkc8qBhzsijqv3qKOuc8G
la9ZdFFUoUJo7541/mzKEZi8omxwo/9H+JykzgnlkVAE7pGTDMPVICCna1BI3nh2/MuIVMM57lFZ
DAB2sBo+4Xu9dRcjg1tXlT7jguEY6WolxswDvhAuf7BzxY5IMoID98jjPMCVBoNQA1ttVpPaJ25Y
FJUWIlyb1A5bVpCFyPoeee2/NmvEU3V01Bt8o2OYH6Sj2QhfMzexGX3i6rjzJ3N19ui/a9nzpNLa
z6GoyFIbIgtFczrRVj/s6AxJbBFLii5a7cTox0+jHanuYDKTdWKEXLrPbtg2oZBs0bpFxau8nzZc
XNYeypDNfHZPzAJJbo6xV+zn6LLbR45zOtBVAPuSDavGUzcES8fcQ5Zdhq7Izi/6NLZj9wO8GFMP
RizP6EuhxlX5dUrRzKhAnfDRGHeTW2Yt8SMJVO5kN7WuQ5ONaKea9Q0q8cO9k/+bcx/L6OqkV/1z
N0F1q9tyg/bjUkm6iza/phDJrQLgNaxpeLoIy2UX3X0+yuXq2Zx3isiGJ8ovq72K4tUY2mIAsABq
H8oKPymGvHG3ho9K1lE045GctDg5oHBDbJ7yuV/zXITLO3L4LkE/XlCiJFi4ROKxO6F8NTJn0QcB
1ozBHJpcixmEjJBXFsl+usuOBtbYhEJS8jJqFr8IlG43WHQ6EzMQnsrOK1S5WbFx37+I8d3OvnZm
VAufduhoYHmLS0HURWoLzscWfjT7Dc4SC0P92lE5DZCIgj+93UiAOXmm5o7KUc1BqNp9qjgnmS4R
kdlSSPzzChhBplW4X9BpB21aPxiPiIGBpI8w3F/x4yeBviN9kt5KZgXpvxKENCsgILI9FqbF1Kd2
CwrdE0UTj3KkjObfRsXnPRv09EKECaVbTfjtPJiQ2wRc81QaNhEECoJook8ZmuPzpos9edb3mV8T
KRXYYth8g0XVcNasFeEpHN+fM778h31igFRnXehfuv1j6ln3ex8eesplSXRztJIRmMZBqMXanphH
pMHxKmjRaeJu1vbTBiTkOA9914Asx4fXwymzcGDZIrDIlR8oDtvKOxFqRGQCOk9q92+iVh0tUKpk
iBqBw1tT/JhGVzL4CDXl5Gvuh4nLFwftV0wpCxwxQURz3BFLNnAD1o28Wa+EZMVfQFXtZX9U5/1l
Gxdj5Bk8Iy/HNb8yYctdWmhojoXvpPkigz/8PpRXlLx3qb/gsZriPvH8aX4/GeFxIhP3C52pIFxx
WdwftRd+hUlY6qMeuraPEViqT6+TGTVzr3FIb58qXHo8jNe9ezxDWZZhl+ORhbbTi+uq3wrjSLoC
QKqWCDhTVyIXm/0rKpnSTMl2XL7S+R5Aa64mUSqbQtGJ0lHcHk9i6TApFSoyygtzALt6YGL9nlSp
73cQ5qUCeBbUxEn6aNA2BLTBCszTSl//8pS8ptiIeAmWB4gQhA9fvs/tK2IzfIOzuYDGJAg4rykG
ADOJc9jlRrY8BN/GFGx/NL2jqPnzkoGSPo/jHl6CET+Ky/IgYHj19O1hFEZvvv2tzDSI7RDEzXyr
I2obr1bOFbv6LOGA79b22xVTwn1cgXcx0e+e4bgFWNrmmEmWx4YkWZ/IbxkAcXpRJRanyysNOryh
h7t7lR9kw+WdSPP8/Qy6omhCtRMmTrX//oCKnbcvd5QstkZF++Yd5/d+BzVQpjwURBLenWS9HBMJ
w5k3oN+uoqoLH5fvQGl1txDgPAwmZz7NwoXSp4qRm9D6ZnbEECHvPULfqzhV0Ok8RSS1NeeMO1Kh
pZlQh1DCEq7pvzwIZeMM9b/VxkrKUxT8futzb80c+PwCQQQuMM7z2COzsTmNWNbM1An1DnpF8bwa
eqZHgdX+ePL4wxTaMle2SxCvJmSSnZkGFl5BuCVz5FeYj/+Exc0vY/QcMjxn1Ho9WCqisR+DkRY1
+s4jd/mj26LJLvfPZP2qJjEvXMqlOA9j+MCm2X6+8PL8K6XR24aV9KNf/Sgj+kdQn5Zij9D47IGa
OxRFQ79a9rSKxXmC4zbUAbinNjh+y6nJPHc0ONfJ30JDB0RzuOHrINQYFQYeh9J4qK6bG4KVRT+s
9ObHKnrofv9uO/nt414z3jfu2jykClThZ+PPmuPXmxc9wb+BpaBcDZvyKeBym8kuOIcIcSEm4TXG
4eTReZteVFMieaN8BlIV+Wpw0uudDYjSeXZmtIV/Lh7H5LSPw+5EcL+0Ogm0uV9Y5KcVQ34n6VjT
L6MR/h5EZwmxaqKkcoDQPJQQ6JvdEkKXX8NXeWuj2lC+kY3iEJH8mkWW8Kjm/9m8ZdFTZDXElAHF
ky8feUAaeynNrKAluv0MiPkHERPGObV5HM6iRkGcOTqrRcmMmWSNjbWJZZppVla0dMlZL6jjFS+T
2T1XpGwgRDyyHeF8MsA++xM0Kyu5CZIxRrCDoc3/OUiNhFktejj+Kh7q2CA9NFTOpJydeLPnxba6
e8XSqBjjzSRKeW9VlXtNUVasojh3Hc3AchGPOi+oVp6xmiK7D+r2cKoff6TfWFToQJYS6yYcFaP3
wJnapPFH7iNKZUsdEJKohkwgWvy1wKh5I4uAjrmaaIxi7T4mHDBjQZDkEXXegEm/A472jSV9fSS7
HQ7168O08Y0mCFZOxZewO+0XRvYcvjyH47tbQjhk8h58tlrmWVrY0l/OXMAnI3ISFMsc/iJYzeiQ
rdFkcMcaddzSWnOq0mEntwPcofTPcW9qohrbPHUdx0oYY+iQbQks6TyXkc6C4JfvuRnUiOfB0Hvq
xm+TXe6cGDhdusbUAtn+1w4p81sFJiD2/7z6UIh9D8GJLqFmHc8YPv/K+fEDzhrDBuogIEaShrco
sapN+KO8JItQHDHC/C3FRG0JCzqwozsNVOe46Hr/cMKTkjTJnHVXoj63knUdWVIGufLVCcjuyG3r
H/ZOci1BTACHGssNLoGzFeSuHRlhgLpTsCqk71o6ZGHTnYIhaDZbWjteoDuxf95yMI42QUKQDIWQ
G++zcDAMMIi60kAs192GMttrecgCmzxPQD0KcswDHdK0D5hq9ubtaA1h7JDAX1043qRJih/TmxyY
QOYc2K3OO0EJESN/oLAE4qtg7K/VmOro/dYq5fTFr3GOAjDrb6dLwwY4yxr/0AG51qsWRIIr9Hnb
l3q/bRrzp9KvIJZfQvO7RZMjhwfPVy9hf5xhk4JXfl+HM7jDJikZI6kj2rfonyk91+Zauc1RqwsX
47N2BnGjnchMO/kUr5Z3QLrriOn47bPcmkR8rzPmP+32GVE3hl/xKSalMyk3BPRNV7iDwKJqxWjS
g07MmFG0bJC5gVvzpI9g5u2bHnV/NLXdTzUzOZPvsVR1M9osBH6dBBYzBrGXiuSgNWCkYEjon8Vu
CUcUepX4nQ+lfErsTkldwGIkPjgtxkv2V5Mu65vRmuPD8lP5jl9vKIkYl+t9uiqWID3DssGupZDQ
+x+BekaW2jRpPPeoMEAY3Guu41mrMZa97L6X0UYANxgk++sZ7uwVdzOeZv/jG1AsrcJdUlyy7AW1
L7L1YXEPBzCWh/zvd1FVP72U3QSGLgZJDQPbGdOsMC4j66gruf1RxrDilEIZR1B0qG0Jokmytc/f
7Tb/EIHCof1l0EX8JWO2L7C2VzvoLwsZwz9XqnBHB/7K2E1UbXD7ffrOo9QjHokKNvuLheT9WqQU
x0Q2uQG7jjq5BAXSmIdAP2g0A4V46cnsjjLc7UF2Ritx2mHwBYDBwkrEB4sb58It4ccAT48B5DoT
GLPeoqw/ael6s8mbaZlYtxHC4lYcjBqfgGBXIfW4N9KSylZqYJnVd9PRs1eHKsvfFBufl8d3hKvr
lpsrsayjJ5AXwEqIT8tb1yvtbxkujpbeWhjgAciKEVO35k7ugUMZ2GmlJqDNvRD+vz6mBIzw+1Rd
FZi9nvW2BshcM9NHRCtrmnLJIGvFDbPOaROG4ELSP1+ULwUoKz5Q103qdrg21gN0LfYYT+3EegZH
xywn4jog1XMHkpYy/VZzYdvbxTBUvHMzTV6iudOjEv85pRp5GdxjjbVRNeD4+3L/EZ+JWr1UZt4a
I2t4OX7N3ZVZS8Foy3f4+XniLVFsw6apvIs0OjQBIMo9X7kDqSDKh3xUw1f5VezKQvV9wJ2s45Uc
4Fv4nWnD1whJH8Zo26y9YqlLrKnQFypAJrh0wkcCGJ82bQ2Szpe/weTsDyuFSfXjxFMS/pBSpOcI
uhhP2h+vELrfvebmWcuMA8A/RfzJxTk+LK2kjZCrktGYkNXhACUpEAp6jMcvDy6QxN5iMlts7cQQ
SlBzkqd1ZGcDY18KyhjqCl7MliR1qUeSYiMLL2EfeifS0fFhDLfYrmx6ganPG3hnlsKZLqJnM22j
umemYQvkPPqqU9V2FZCPHmBg3204/j4b8646pUCn4BnE2mBTlYQ2C2p+WzNTTG8KHcwutRiHhKV9
rZHB3Ci+K3cOjOKgvp3jQgjgGZfCILUsrbBA0bWcoWAQuzi643eM/vdLwvQ/+jJyvJLTPrB6f9St
PoRsuG/ASCbdYiyximWGVrHhdCh7Yv2D5RHkiOUCJQRB41GfDtdg1fLjjIDpDw+JJFr4mS0z0tZB
fO3Wyx7xh6uAd18hATqld5OiTRLFrvVo3SXczByYUWmMwdzusOZeHeDPMF08aR1aNi8SCNaCMVou
9zyVoxBSG3BKcZRCdu6zYAgouAAJeUVP7YMbFmy+qWO5qysfLD5jwa6B+tgISOQAmT8aXXSzT2Ij
QXBzhjamOAupVkhF3Im6UtdkoRFLznewV55OTEAXfKbfpqTNs9mG9ftMZq+9POYzeByZKJRchQ7W
aPvAWN5FOoDTJs6Ce2RrU99ZxtMfJWmv7vtr+me4KelGCBYJtf9MnJQSc4hwJcCWA+xZ+Y84FhLr
CWkhJWRCDwfdHs5Ujj6hIIHgo8+pUvMSMAzOme/5wS/JQ7pHYiEqWysDvSk7H0LGT7rwWaK2kodS
FHy5As+q3ZnqyxeehLB2Pl2Hkww+NXPHhJJrWVGwQHdz0faSXvEsOsOkgfIanyZiO4asq8hDgbpZ
UR35lQ8qovotGCA1V7wptXtUyLfyTUkO7A3orMTl9+T9InFWwMi91hYSwRuggSBRiX8gqLbIw3wT
cyZI+pYN/rganVcMavei309o58KVAv+VmSCAQUx3LQgikvZyZlum13FAJJKWD4OQV/n5Jk9mtso+
XX18XRqF6l6ypR2sO3GfQ7u82sIE1gQVDerYP91hAHjlZkTbcfFc62zi/o6AM7ghGEA+GBo4lxtu
cZuTCKHF9gcaL8GCs0H6RAvWrFKBcZ6y+Pfk3ukonZKabAasLI3UMNvWal+Vo2vTxBBDgLFaZYRC
bo6ByfXRb9oWD2+F89edcZD5XuMUCRB8fmTi4g5txMrBkykRDMbU8McoGc+c7d5QAKpFjjm6W4H7
bF1xBYhaGLY23RxaXvyPr8abSffA/KLfReMcmbRhS3s7Jt1/EPNP/Ifm/jPHIzQ+VveO72vc6gNk
zl56+r5PQTJAmoxdB6SuheXoVWQuFqpNtGeo1Aq1J0ltXP68BFtqZgeR980Mbm/Bo1Wm9dfa0vGl
hR/lfbdn84D55o5UAa1UKZMHmeRcVX7nprLR9g8l6X7A2ovkKXCHNo5UBdBVHAzh4oRnJ/QB4HlZ
rs4bPuxJ7Jfe6yAJcaM6aJzwFRCaAwRazBcXycjPQi4ESxd55roZVx1ljcnz47KjJFW5Q5B2gj0a
I45+/8qdyzAN/6ZQmh7ItrFizX8UOhlngGqXa7uIt/KtmNeOaZx6LQaDYXVNBO96satOymsMuoof
VOB+NpY9aZBnEGW1nK2z/gJCZlk0BCEghFqTGEfbFCbLvrURwTE54XTt7Il/Y2KwaJgR2wiUCMUg
2qzz7XD5ZStWTLebz1o0rxQHScKdfms6nl62K5ygYL6LRD42Psx5fbAlU6SCtsy6OBrS8qoI0ONI
Y+gsK2hgDVoMA9iru6xBGIAnPe4FCsAhfTwEMdhA68tq9X8i03BqMfTvU90b5QANr7+oN7gdaOcQ
xHdbiY4Z3H5ss3860Av9/LecR9VtPTuV15hGkp8RB2BoyIpWk8Rx6+oJ18GL9AdWv/ekey0FlVcP
OcKDzW6NKnCxi9EVARF6w5heM/GqwPA6rXHTPPoiHz9SVKohnumulyDrUVdH/HK2vJuB/HbV4G8M
PCmaPLw3WKHj7D37hql2yL6aGBTY7i1q5EG0mqeZbk9YUkZ465FRjZxhg6uUZeyS+RBRac4IZX0e
sqLDK1XcMUsCUAIdde+IdYIFpXPTo7kouvw0k381bcKn538tU/1egh6AQydJJYD8G0dytS31+Z0c
nL6hhv2kojsqFymQkVENYb4AIuJU4sQCQqJFIOKF42Of7evILfcTLZywEQy5XLs/SuVFFTPGoQxl
jmeTbea6EVRH+x8qgq+NtdGZwyz11shBRMQ83n1cNaQ1jOSv9pKxcus0F+xagUfBwV1Y7N8jF1sc
rtoQ+xLsmCoZvIg7iYDBio5LrnUzk/maBUPo8nLH7Mhu6w5AhZFU9rxUrsR26pvV05FCmuaeOysI
wpBzPr2Io37/j9HA0lzLUV/czX3fraQZZ+EVz8oCYh+OGvp333xuk6eIOCqq706y0g9+o6GRGDpl
bBgcIbLvM3Gy+diFUlCY6s9KwvOHSqKC4m6kR/SLv8cL/R1n9lhDkdYdS1pwLPwIVX9ACp177z9p
duQ6kEA9c7LqpUbTazUq3sOL72PzwbknGSMljDEp4xgsACG8RwBiPDLs75tvUKfAYtF/0micpsHg
+QLmMv4ODX+5VBQ6ATVmgWoBvZCorYutUl0irMAAXCCGYs0fGAllsURPjgdx05TbDzcpnY3XrOhw
qX024NLr1ipOuPpQB7SIGd/iuAsc45jR/ZY1XLON9WTzf8TK61cD/2WaF9C2+uo8B5EFaRMkvuSZ
ORG+hxroT2RZktaUYopJLhsg0IdI/viIwtaskXPX3+RF2VNrdX3P6Zb9sQryD8SFLRCp+iYfhC7P
QyK9O+3hlFtdRUcit3Le1vZ2stOtYpGibE/9rfaEzJCpTppqBmSXaIPPr474RjrujtuKhmwe8NOd
XQd+T0/lWbb75ZzEek7yNxT8XJ0JkzMTWeD2OoUbrUk0m3IBZrh8A+D4YxhaNsHOF/zqRcnmglXc
13/CA+NKE1gjYFqMcQeNM82NskaGPamU/fkxIWq8z1Bp4Xo6KH4ba9Ddhy1sNSTrVcj49tCyeYQt
C6lwbjoW7QozBEt4wqEPfDcuFvS5701a4FOleE+VGBsw6oaQsXoa3scasI2sc4H62XUjJDlqBV5C
AbL3XTxk/FJmAcMeb5odwq9+jMildVOSXW2A4CjO4b7h/o+d5a/uYuKpJ72cqbu0S903G1JD25RV
JePrFeSWBXW43swBizalt6d29OIgnzhZCVSHKLwUj5HyJD1ba54zmCMFQcvxkeXSar8WkfQRENAM
OgLAf4cR5bp8fUNYxlXpzUqMzqOci+Zxy/c1MZ9ZqVTOSvOYKUpEwq5J5i5InLFU91JZ1Ctk5TS2
+Gh7dCYRmdkWpJIm1RulW1HW9+SPma+mUVmsSIv3dLamdOy/RDjPA+tnwCcAoaJkskeWTYPVuc+B
+Uj/gFDidQinbci5tnQ2nyMA+xPXG7tfzqp/mpC6tGJXC1fvfC/r0C/+Eg1gbAO8NKenca3V8nHU
GmOfLuSQe+EF7ZxQjdNmAmOip64eui1ASSdpB5AaKA6y2HW/s7hmud+QiK57k2A0v9kQmiqfMMI9
bc8LcwIXCkH31Sy21FlN4/xxG1rC9Vu5F31fhuGmtiC1kNmMCJuRB749osI6oONL1rnJlQ1uZDRu
sNDoQO5oCD1l3YrC2RpK6Otu1pk2sWIzRYrnDNk+zsxQLwmB7ZG3h/jCY7gp4BOzu7BUROlaBis5
kuxlEzhSEqWz8cavn0HGDdNcbCqj+PQjGZhXHayGlymYI0pbjKe1sFwysS59ELnmQG1o7D2KAICj
OrJU3xe4U7oAvGduj3wV3w79icb1XSIblOQrjYHxyAPtkiDJTA+aRRB0AxYFhEsgpSPR8gV6+Vmx
Cc0LuIiK5VxZjqmSiWW7AugxbaQkkoe+eXNcyMz8vCkTbMFnwSZzMKs2QeDnMYmBYnTsBD/oa8Gy
ZYeN+T/CuDMxQ+5sssqiLjBrGFD1t/NsjrXCHWSLbsDuvjCu5bnYVAQDyJ4QsaoZaoOKJx60uDhu
FbOniVH8wRkkeXtQSpqVJCkwjd6LUS0TxCKQsmStjrWLiIKa4VqhPO1S8iCC5tkCVNFNCTRWbei/
9k7wx6E9kfmjx5yN0N7UQtdOfaG3tgzWUMurN1QRK0dSDKintMUpKHCfrtEwZsfarYZ46Z3IO3kp
FINKcyKBLMkQUqy+ql8tsCClgsjiJXuCdTfR7bBBoPcelEtg49AeaccKLBMfqLkow/p4HTeVRHC4
dG857aPt8TtpozFcbkirvrFwM1Kgs6NShJYS4lfK7BfGO5iiHM6ECe18+zVxinJhDIdxF47F7eLv
yEplL1yO2WN8ZBLCQiu3Yl9lOPMdVF2i8lpVdblfSlHhNQ/CmquuZeXBf8RXT/a95W1OqL31RbBN
gaRI3ffvNGhKKTetdtFtHIyJCVJaqUEar0g2TKZ/IEFellibtzCYkgT5JgRnNxHj3XzvOwEaoaqu
32DKxiQlcq57J/MljuC964umPIM5QW90Z5wRbx5crvYz+3RKI4PHwHu6MuzPZwEyjpsgldmAShcd
pgCrK+uf4ye2WGXhAVQeq2AXAnvvvYIKseaUIwgXuEZJhf6FbBo0+V54yEGqbhFpc8ggD6Y5PDzs
Os8jOj64o2W9U0yOKyTHfCB8pYKf8pc/6+M6T7o/8AQj0K7YMvYVryKYw+EQjbdLnkFlYsCKh1jx
RNk/9vLACY3TVTBiEUyRs1Uyz6WhUWYjYZRum0sC919MrBVseNB32Scc3C+acC5d+JDYD0D1BFKi
KRrFDUW568j/i/LtoVCNka8ls6r8+VNtT+TJ9F5jI2+zK8EOWEFm7UDYx1gDTIvVT1rySSwr0/dz
/+k5ELKsvwp9p8/yqpyaaN8rpOm9TmDj/zA8YsgLsVrNFM0vxvC0rLfzDokVD/ni24rJ/+86eTPU
E2gcvpKMgppQVZ9MFThb1+5AHeBgBszo5k93F8aa4BAq3oASamcbCv2bsbHNJFd6eiDwbdmlD4Al
W2W3OWS8aDu6tvtRk2cLX+SVLHZ/J4QyjJNHjPsFzKqX8vk0FlE+ZIRpvX+HoP+AnxGIUy0bAhlM
GR2z14UICah+aIlk5juM+o+QkXy39XJtw+g+7eTAwTHbXkGpim9c7AAxl2bIVmV7/VKxGZrCwojj
v+Z+sOI+A6kRwK9SvRYq4ixrsmqd5UPCmMKSUdcQNZZkgmdgnhBhx3jh4tWSp7H9pnt9LqEFF/rn
vqSu4i1hJOLkWK+kNEPVJbQT3CMnw/0KSdpkH6lyLgaHLLMV0+Tb0jNukSHsVntsy/Va7yXdzQR7
pJgixTmtsC6h9A/j88mZDj8O+F/23RzHXRYvVCgE9bNcXnDh9EZZ30MFaNGQe9xIcAn+R/eXjP9F
KewBSBTmz0YWhbLokm/IGWly4oSxVlija8HqA7ksESTUgGLwoO2TJ/mbN0YvpC0lQIpouaPd4M24
N9rCItnCz3nqFP5C15UuBq1CioopAX5f+ALWOGIGfHlYQxodgVBkDgUrFduzhFHA8ljgMwMKMlpM
0meeq9Md1Dfg4LTJSutJMTfQYxcXtVT9sEpOYiuxxSg1cwkmHpFhtc09u4O+ZvEybXP/rMhlvGXn
w7mCuPYvwLs2oS5VZlfSO81acRU9DSGH7GWFhDvP+GKJVmDBtU1+jldOtMMH3wYcQtwB1aj6ieqN
odJpVvqEKeAOxu4TX7tujAVoKVoc1kDqLaaLW86AOwvO12XHK+csXdRjByzGyhQ8mJ+KqCvSlTH+
jyykbD0EpT+D8ILf74LHvtbTdGNBu8xa4sEdSNsOG+fYLg2NKDwg+l/FFJmA6lmILFjGkVL0ivvH
kRqRQyZYmTgHZBTRcWSqQW6KDwZR+c4AIwvYMnBf/TVxAqYtHDmSIh3V/ZtmchtxMaIwPCQM9a/f
hNaAOMk0g0PRnqao4NWvwGJt/drLR8NIgL46Cmt4McAcZeIvG9ztadxmcuNYFymhpjoBThnsFq5s
MgHIkgVci1tGDQQilyC3YBe0mcXBmhCfrqPlO4Sk7wMBdJb+/zl/QNc6+44aEgzruZ1QwbIwGbvL
1OXr4oYoL80Vev4v2RWSlIQuL5ukgy9od3EG6PQYdg3NPUiJxwU9P6NO4wDVhq6t1QZBNwlFSssC
/LJXub8hBHSGb04L8pFu0wwFCyXATwyDyMW8tXLAksevv0kN122rjk6kgTjOXFQ6hWbh3tVBoGEl
9SItu80v+bxhSmKCXWU4h2KcsDQYA85YTyVDSWuCwHi3mhQwL4T00z38qA1bRkMuNMsuriRlz+Q/
cVCJmexNwIm9adGbaA48Okdxs8zlhvd4QM7vmrifIGFVu5kloDRGo5/a3OyI0iKyojkcYigsnXKb
rwV0k6EecklKpfN3RiXKqIQrruW8VR3T+3g9zaUrP4LBc6zNP/gBVEtdkRU6eSm1zw5Hk3xr8iZq
I3LRDWuJdmkqS0cpsxd3p6chDN7q+Tl0Aim20MSk+DCx++x1TAaEXCR1VrMoWRKMrCtw6OeXsBcu
ZU2Mf75zIkZFmuYk0v6YIKH7ljR6hvtNr1Hy5Q8gip156FsoVHnEXl/FFrVWoV64XKvrDvn3glXg
rQyZOpXWCEXPt6SqSxwSRqlQX+XjNfI2kDAOVQSj+AiPA5++bVxhiMVIQBbMTd3kA2i9n3QqzVb+
S+GyWRCD9Zj+S4iw2twQb6bjoWYMdkSQq/QERj1nuHfRbXThbsCGbLZVgA7KsJ2AdBNNvSksO7SR
kXuNA+qgH7h2whCmUk7v5dLcmuBdjCCdkMxa3Gipa83LCDB3P84/INDJMR0gjRzEfKioR3Tghf+U
KiZCEMWX/XF9OuXVZWPH/X14MqfI/uYOk2uT7WX9D8NZWrr3PdXL85jkgGfKr3wEGri5/RBNreWX
T95d81R2jdXihzbzxO5DadwMZ2+ebHgzapbznnypdZ8rmPCjyltFZGUQyZ24fdy1RtRbxc9pUyB1
8dxMP9hxY7pl5OpHSESrA9AHhxog3wH554ca8WmuNRrT7xuluHKbh2Y8yYGg1zbFJ12TPQRypBtJ
yaikNUw5Pd78WTXVNyMOLHQmHahODzAtgjkcAE3RYjFd5prcQp9QtqIMggCQHntr9vrSYGq9/X3O
3R94fUycXPrCnxqxgM2WLM3lFt9Hvqi/QwSKR+JDWYo4nqcVfdc2kbShYUTyq0OjITwIl8siDzes
V2HEh0ZqLtKs3K2VrDhx0PUAKQY+vZWIaRfxRfLpGlKp7AP3Ll73R0KLvhCdY6b5rmiWMdu1dry6
gjoATn4LCvbhbKdPl7rxPUexaW8zB3tN+PNsffjoq3KYoVkQjKtOdoAOC752LGtz9tYx8j8NOcEW
kRnAWXVMZAU6QepO8Q41kO8nCnmSiqBQd0pE8u1GK/9jkq8NOCIQ7kbQlob0CEBTOixzYus0dsMN
uMTHIIGO7gmSlKNLRpG6sYnIzX41/K8grRokCD9qoawcXPOjya8fFN1qKiGhoYkz32BGWvdvcvXX
8cnRhoQdRgm9X42VX6HNc/WLgHzh7Z73zS4Ve6wrp3pg5yC/QqqlmM859SIuEbuB/A0OnoFO6m1D
MjokeisStC3e6Co64wv8R+Yk0ZSChGPJihb/nLKKExo4NvZVK5Wl/m09CiRXtjJyDaSNLZr1A2pb
tGftaByFLgJDPtW2AhPFIHGKZsrOr1ACq7oZwsC7rBkqZtyBu0Ga+eBv4ePEduBAJItfUke9OW18
jqVw7aV4KZ3ZTyulncqKtb/inCRuZiIjQw37zZ4YatTI3KIzsWkdKASW8TJPEkm3sAnyNGWhO9b5
hIrgBUR92oW6xhkc309+Cehq4oBnlw16N6Cr3jaLr0HoUPjYM5w1y0Ab/N2wK6ZqhwsbRpjUdzz5
VYVnZHUIgeUyqpBhLcGI8w1dwiCBGCk48SCS8Vsa3FmNkL/KJCQp+c89OsQyLxxtBfSkzC5fVsfM
vT2/sT5uexE89q8Y9j9UBWO5B+PivlmzGX1JP485kGbk5uHDiyhr+hlgHkZFHOa8ABzsUiOWz/Oh
ftNHnU4rzWbq5/0Tua6zGixAoHDJP4yiv1uVv+W5eUeBgxgXDazSuv3GiYB8S5rXJGQm0j16UNp5
MIZ3kkaU4yZ+AD5t7/spPM+s2lxelgzmG3dZ2hQhb7QZ7KVH/HwWbhCYLLZbY6ef/PPb5SmdLmn9
+ciGlA8eRA/JLjQ1ZbrN0+qxjfOeNLopfMazPCwyLFy5Ha8Trf20w9vElRKGUFOfxmG8bhgncy2m
utmuQ5rrWA9FQF/uWZhGqEJpSi1ce5EgjKhQ9n5ITy8Q3UUrtNcIP+epghV1gg/EiVTjbxpKAkva
s8m8nDe2tyQ8GQMu21iW7AoRDBWDfcE54T97Oc/SdOsIR8+8GwRFKW9Wys8UZVJKjqC2mL5NU7kx
rGoV5i/TFWcgKHmqc3yW8+TI89GdUwyKN7pmYoynfhtt8WXrygStPnPThvMYPDs2Hl3TyyefNPN+
1RBW4YUmbochuzmz0Nz9hUvG92kCqa5CqHmmTur7xppBkrJOokXKmbYnWC5W1Jd1Yaah4VAKyzl6
/ltx7aeAH3cJYpKnoTp7QwZ7cz5JZOy8rIx38K+VzXoxIlyQ1ZpHUbgzvbEhDKuNqbPRxc6Z5EQl
ti/BecPoi9mIYrwPJcDHZB9MY7FAP87HJuhK+VyjRF3H0R44reVi2JrUQF9592oHqqi6QXA9t9sv
E5Ha4lnb7/ZDAKQYITZuvpP8Hf7ET4zv/E2qQN6Xdn1LeSk45lSLHkk1wCgUHIjiuxroMQH3DpfB
H3SzMkP/TQ0QIjzAFjT8LVgvMMo82GFpWhRh3p6F8947cXeafiLH0zjUNELKO99R/TiFDU+z25GT
ZT+5jMGekXXVkbW8uhPeqsg8D6CbW4EhhGfAIQctFczXvTCJaiJE7QBCG4S8trfQ4MTtm/WNSGD4
DlwC6lYCxgwoDc2D5A/uQeBuYWI6PXVl6E/QwRT49seagO+Roujh4w3EX7z487kgb4+enSMxI5uB
/WMCteoLoWnb2U8MNA5YYl1qyiVVgnJbTAIjKkmu1/eE6fTQnCrKlbMb9AYoI5K2lUOMhr55bgI0
+/xUoye/8/isDPuVaRsTaRogTaoS2pRyPNq6iPRuxNo79ftQ2pTNieGQCe7TsVV3bH9VsMzxswGv
a8QBlttpbXdcoA+SyNTJlcRrtah5Vwxck3IQHR0VXjlTOl+1smY9yku9I1z2ZLX29mIsO1m4EvGJ
StcEmltf4A4jGh9/uX18xgyXRXuiTiGTjKWR0kle21VIh+yu6LdsmYkPCMFvDBRLAWUNlwRBH6cE
KuuPpwfwdCfAsA9agPbA4TLsLmT7vvWMHTDfMROAwEHKj/XUr44DSsmadnmnIbVhK/0zffzmUJcM
H9K8rwEz8BGRqZqyamq5liGnY/ehDehi3VgCerarpbyOw0o9zhtvh8vtF05kE0W4L8b0GakfYB1e
W3W32INp+clu4Sil8zgzwXwyxExTqOcVRZUshKFSTHYjnxALPnZNhiXv6aDyna0hko84eSTsmYyf
WVe8eWnZmUTl8oeXmX6D2GPOPLOf8XMG/g/IKwKhFOjZgS96xWuZgc+TUHCeCUx9AgC6Ez7LuLob
HxAwqTzBvjF5sIQf2J7AynudLqFU9fK91LYE8Q0QpDCkrGP4rSfbzzScZQzGDpNtmzdJlIKwDHiV
eXDqUnaMgGl2pst9WlfVFHCOIcoaItSeBGG2O4ymHFnsirZLzMiTdMiI5X0wqYfhD3sgzVL6gnsD
nWhLMtF2hpBcmbtZxFXG0RN3HzvKC1h4bICSH9v/sdo/ijQFZKG4F4CVOgetVYPmjJ32RliJ1WAo
jLjulmUn9Hsl/LUqdPEx6Z84wUTCICiefUOlEt8JT3cKva4CfwFuzLzZr/XPYIqDe+d2EtdUl/CT
Y2w3vqu42MPFdgf5XBSKleLdLeYY08vRrQadndOf8hVJxQgrRZAHK19QMPLnA1G/dPjhH3iyqHKx
nasC0VJYBV6Rf5L3QiZhgI8kN7XZr2FBsIWBF4LKJ75V6egksPZHR6lBuxSAIBViJsk4t4YMYDGy
8oVwSEP5e4lHwtbKUX9RdnC1uZhVmTeR2x8czLtGkx4k1UhD4aXe9bzN9SoSl7YIR0ei+RZl5Tfc
GNvAgEAA+C1TNlpnWcxyLD6Ic9Kh0Sh4IZf/Awdub58S9dE2TFWOJ/I6RqCVOT0QFFpNwW6YHs9z
RQHArT5Xp4ILx4qWYP+iEfZk0eeB6eIqIypGoaf44KWLVyIVdHyZ+MLGpR14xdXiAL28m+uxbZEb
XwXl3ZCmi58OiaX/4Ds0+k7x637V5PC/MvoM5wJN7gGW5wr9tOdT2kW0VLR+ocln36nxqf/r1I80
F28Cj+gEy0Eqc8/AXrJKfa8pRiiVbOXlD8tKIzpXIIcsKLlVcbeDZn1uakL4yZPLmMdZFIRNu4S5
8L1rUhl6lpaTcHFpuM8yHGK0xhPW7TKfUH9NHtLYJtFNfwxvGdly5B0OUgA39qlmwZM99Y3OPN0k
6O+TXwM9EG1SF7uCyL0VNejFovzdRYzuBFKr4NSbL3TFqZq9H3vUdcXUuhDVaooqkWkg7QacUp2T
8niu780Mw6nw6AKjr767qKXseyZ40+JjLaPW2QJXfcnJlfw5dXaf8n7hL8CGdcAaZt0BsuQIfYkP
t4cbnyDR2qhjMJy9goc+/Q/TkhNKM2j5P435e3iihhwJQt5CNJ2klZ79eoMncMcmP9YilPeZywO6
30a21oACLM0GUpRQUSy6A5MS7YAOzOhaipq3kHkuWLNhp8RRmZVkaf5EAMb/08ia9mLV2qSsyjV9
XNJGA6iE9BybkH9K6D6xV1QM23xD+ffPEJfQtxrI4vUmAjw2TQKZXHgpf3PiiZLF3KuWtY8K8iNQ
9cwjou300Z6N7KwekKJD33VfdqUvY8bqdHsl2YV3BjSJgKsg6tn8okPZEydH8sM/QCk7jbqwGsd8
X8E6fHGZ53O1ygq3wY4iM/T6Tqv4Z+oKa7ETfEFci2viHBoCky3Wlw7Qu4G3L3tDD1X8JVhrxqaz
+oLSIoUFqGwYbI6b7iH/XgGmeg+cmt1JpbZa8OQb6Fgz4iRkFNIZRl+NhpM7DcXrowiICN1nfC9h
3pqqkPlUxqLUFvBwvQHXoBOrXj+dhgYIup1ABlfXy9soweFmBqqhk5wjd/G/icPikrDC5uCUIU7k
6yF5zHG2/ifrJyBRL2YiPf3n/uwXGTmANKDvZOii6Md6UdOPbehBLMagq/D/yFiUqNhHKIsMVHG2
lhalX45e6VCI/ryIv5gl6GO5QT2aWZvUTZGLzyZKmcMKvP60L/GidTGQ/RwqhFf5TgTVAK61lExb
+8AevuMqXjjF4Q9KV6fMUm3ZpISNjifOnLu4tt0bzyMdld+yhtfqSvfq6KDIGiNzyPuykzK6nsbi
poKYWiF+Jh3YZ9ra/U+B1pMC+TPGh7gNI5Mb8aa2CFe7bA21dQ3yqF9z1Yojug3LcHhYklgOPdNn
s26gZjyWXXorKaHGdhn05LA8L1tgBE7qBwLZepgIaujB4TLOrYgzHaWHRQtxLnacX7G2zB4tANyK
aP1Yyv3uj0groQ6vc/Rx2hse6XCK7y/AzzrmhHMbA4RTCfPn1m23zVP05Acnqybs2K/WbdmWoCB6
P2dIFYL7oyezhBQO1RygNzZ2uVUGAcrm44R3fbs3xt9HHbjxZdz0bgWW8z6xJua12+YdDNbs3wUg
ayOQhfP2hNZ53T+U6YTOgIRF9k7QnQb9a1elvTnbdwq38BvnocbImRjcM41tgzaAK2H7ytBRKC/u
ANpIhP3sKNV981wA2TK0XSUjSuAiA0q824EhFfTA5/R2H7wtarB3nndzadKN2EppTCINjmA7FKLu
RQdDx12Fw98TKbV/VQTc86CiainIwz1TVl4LQTrjiy1QjpENjobEPN4/KDbUs6tiGxtoaEFi7uht
7lqBYTZt30Gw7pi835JvOaoJd06NzyRAqsc/Z/sFWb3rZhVCmUaq5wvnpXK4nHZxcqckECw1LwJe
VnaIl+v2wF9QgOiN3cBCuXdhh21vVYAilBol13fQxkDl5TL0ACFax2wiaaM7Vkewo5PjgOuuymBo
R2aCnzIQc0eLr4KM0RJfOVWzbAkee63igxRLZujjt1LM2u61c8SFwae0Esk7qG9nlsgCbhzSSQPv
wtcUbIiRcVNqf8C1sQPBZKUvInwV6L8NWoS5QtrCyZdCjcOQ50hEnWDp7ipAVZVf1eobWEz4ZO9A
7iJWZhqQm6hPD+CCdE4TNs4SvqLW5bf5/ppD5HfKYAep4NjWwtqKASQNpbwF9At8Imu6Hrgu0WjI
eNYyQeE9EZ5d52xjUf5VzIrxjJZ88ODrRgUErTpw3K86LL0T/Dl+8Ypms6rDBDcgnzxjUUAOm2tG
xlCMeWHoyeVO7/8PZop0lnvCqVRUz6EMwLSe08qknssLIuB45V/AT9CGXiJCZQvGpQt2++ZGT7xI
rvqWFNMZKKVN4kE/L04/pbdlLS7kFDU8r4bzBEXvS/FmBYBbTySMCj6L0vIFPENaOhpQeCGhNuVD
GGBU5zKCHvvj4/iW2eLzAJOzkvTSJDzJZh8y/b7Gd7KwaqvxBsfzD99B5/WHc2iAn1s32MIw7Ze8
hPEDrPT8XgtYrilfPZc6TV4N4Z6nVHV6U1gprD5VaCHBxK5MeoWDJRwTBg1tt9vSjCcmZxuej9Lc
XR06Mz4Mf1V56Z1W5HsOrMjvaAh+Byb6KNa4SgCJs3xJNF81lMLRGDrEpmH82O8eceh2x0Uf1KD0
KS2oeFjn+nxM/Lsv2TITYsUAIMChwOUx7VqR9n+wLy19jPvh0FderhkvKtPCKkWo9rhX23Qk6WCj
t2sG1A6F7T2JpxtZn9GO5StPaUdbJGHLZtRqss9pCpgGRc5mScGD8NasMln8fZ14eXnyxEmT4d4i
ARXU0iyTKqPBKMlmbzNsXXP+007/lW3EzxME9ePtm7fEaZBoPUFbQExuV/KZruodFYwp/u3G8XIL
2lXHd/j6UPg894oHUANxPceIujniYytaYqxgR1NUB2SlafbdxgNjIlIeo1d3YVEKcPQC4xfYary+
TxIA5o1xHiWvXhhALrFT+CvzHgmqv06a6ala3VfY5gKln3bLkX15zcpSFsL14quaepPxth6qaSmC
QDhQmBZ59H7RnRIcgEHHfyswOxhWhdZiwDtR6dogFcCpfAyudOJwIIQpknWAlPK64H8XCop22LcD
rCVWqU/qWNC7mFx2fGm4zebUYYrnlTCI5/5+n8iHH4bwEuXNqSFr4yl/vG+3xp5R6k11EHF6CVwp
MYc10YeLbVG06Deqxanv5B8Enn1hiDS7dPK2Mtvfxqd3MfShmmJCYe/Z/E1s58fl090duVCxNRjl
20mJ7VxzHQAqXWci1iQjEQ/QsU0PkEIS19b8lNNR74P5/yjqloU2hUAZhVCMz3ZRUzcULJUPlP21
cfF8EZ/Bo9hSsRVGVa5bl4i27cUQYekB64qIT/3cWIPrKalBDOZmb2qlTF0Ci2R/jLZbsAcMJqDK
5JiHxxFz6Wqri1BGKOG58wMcQmwOJHPEiuKIwE78f1tlLfHiGPbUR/sewEdZt2rVTazYVUbo6hdc
o2/7VH2zWe6N+Ed3C185YDh96BK4sTiHCeV5vKoYMdfulkeRQW+i7KtGyCtunAImTlVw6Gomkye1
iUR0Mk11Z8zE9yDzh2lwrCl7j6B/IbGBquuqlDHtUUgLAEayusvpZJkjkO6Z/fZUxusyNDVKBJ+E
H6n6BD3wYFCqzV8SKMOiZ7A94kd+OFD1t0D7JQ+wm/PhrEUXo9Ez0LrHVPIIHFzPLbslk9RGynLA
KX355cAhF7SIOjRhC1QoMDfxsbnZ5+Yt3lpa/L0BkdZUncULB6en3qclcalJwNOkGFZdib3jcScT
8Sor3ZqUkBs1TxuZx34ca3yjuzBt7YoSXJN8ob1vy5RJfchC6+R3onAY0RA/o7RFowKopy9Vsm5A
naY31h8SYO1Qt6krLoKEi8Z50ZbQJbUrylBpAGLRhlBh5iiHxKF34SkNdS6cGrBHmaaTQCXiyANo
o0sSzJRE5Ih4gq4TNuPIHzymyD89nfRj/UIuMYEzfxd+UC/sV4/YBtvsMasY+OSfFpbSp49nk35e
KBQ0ZOoi9Ebv1r63X6fitvTmtr3v4t+F2r0bJ6YBf9tulowd2u3hDvw5zFHJDS6p2IfDmfsesgds
gFzg1A8GMNk55Ikz9cAFG1yxqILZjCueBfNpV1rdxZd/wLlMfI0sFS5oWGkqJ//IysaR0crkHS4n
x8blMpkvbWwD+jX1fVeplBQXunyjiNOhR/Zw1vbGE8/T4if7QUCx26Fytx0SeFr3htzvYanPFVLm
IOIm2Kr6NIERZRu8sLwGH/dkhZoS/CnmL456+Pk8MXWPPv+du2Ojt3kvFwjwI5i6k3N8y4YSbckh
OjyJAM3MnN+r6MXf9EzxRtDbYkeeMY3beUJuFxyBuzVzEDGyso3IfuQ4U/Dp4jCbDLpftBm3bkR+
mBNQ7rjHWLdP0J1PJQAbk3fBngWQf259OUfsjzaAXpPf/KYCGgtUr5K2KLK0cCS9O+pOr0dZ8f9u
YwguhmP+4l/dynbq5JscVMf01ANxXdJgan8YlHd1INfqmye08hWMJHlCqK766d/HD805e3KCHyw0
cXnxODHZw0HQb/5Ou73s4YEAyNJf/FdkkrjgKYWNgPC0TJb8x37+0ktxMkTY6dPoNddAgOhN3SID
elfcrhP4EGUDWP7GFq7Hqn84vLoGEubyxqM4jTrv9Z+pO7FfWn5RUF8rH/QgqIV9qyf2/spSl3pH
P95iL9nN15EgBB9j6qywUNBYE8xRwDHRiFpJDwiSwZ9SWYc+Ll5K06hFfZUfG7ND8WALwFdkeegf
6zIvUj+mT7QbQXXuD+ZuC03uY9M0LwjBWYZAm0DZIHu9JYJ8eFIqEsfq9TyKRfUUHx0CNWjlRyF9
d25f2iDG6Oto7kAV1XgUtBRiViFkphiM1aBLf2Aix8lfWJqWgaC3OtTcSG3ipuiOScZm9ooHZIHN
Hp4j96cDtjfW2qDVHUXAFjDTkL1MmuMYrwFcct2X+m6G77aB2x/nOTb40TgFqfHbEqqBwUy3oQlj
0gab1qW0X45zipEZUeEhlxWJHwvhCB89m4smMplVcPqlJ8+FzGhlZL+9Ppv1JRFTDsOSYKQkeBXI
qJkgwAVaGfvVlrpS1ObkUhY5FiJQDHqL8XV+JkXLZ4+/E6OXJ2mqpHsGE2eymzH6KjSMl67amh0m
bckzTJjnkXXUA1eku+e/Smh2LYski6xczTUXtbHmdsBw20yVTof19XCfXDS7KTVhxlBBqmc31XqN
HsHJjTrU+ptzGC4WFW5vAU56IzQt5rpWUwt39E88Z+CZgc1Q47puhH70u3+WoZEIXHG3AsIGlcRJ
QzhOjUpqz+G6JaOUTgq/4WNt4pd3zaKpw3NqVKIRxV9+2chA53Q/B/TfExmx4jw7bRQ4sPDS+h0R
MAR2CBqzrUsK1gTAB2+hOW7hKoYY4FTvzDOGPPQiymVFeTtrvNEXhzyz9WUzQ1hLGBT8r/EhHx1k
+JrWGvW515Kxm9cfy7FK+NP55ooQGuZxa0gbPsFxLKZ75G4AEMvzesonLQzkwEd89oEVy6M94auC
v/R4J5g/hzYvtVDQ3lj13g0Qph2xSzDO5hM92zevbtzeVd65TCxlYYIZsdBge1aEM+JxTA5k8TLT
8+wD4yl8VHz7m+pl5+dygvLMRD/0S9mzEaOHvHHMmgUoOTwEx4kwNiQFlWYaC0z+MKYFTavDGe1p
H3UJZYxJeVu1JTLSo1dYtIIJzFF8zo+hhmXiQpGV5MVWWaUhYa1RX9KdWzBMJnWktaFTr67zuJO+
NcyFva/585FMIWt88+K9j8sbyWuUxvB58hTqs63FK8N94Sp5X1ClmGCxJQrlhw4tII/NsJJM5jFN
LeVtS2eibtkDevxhBf14ARj8WAOD3evedDEZFhlmnrOoey9gE+Vr7vSOxtTp8IjEeuiw0stVyI71
DdOVkfm/r02kw9RXukiVLAeCdUu0vPpIIJQeHivHpDfGkWKVA1Kefq4Wl82JR5fyhtMWO4VXiFnY
V1ijgPW8V8R3jji/CyXoQ0ik1QlkHGEZ3emisLKja29PeMa3OcXU9LGDRMwi2QDNnaDtzRurFUOt
wKLzcpo+vmJpLO8URaZG2gX8ObVpxChoPFb3f4TNosSygqsddVlO1fj1V1HieTFwSPCngU9jJPPN
imao1E6l8AeYAzPC1KQIm5MWrihQuKoEnKZS9ELLqq7msrFDa+zDZjX6WVyx6b2IALG/LZ0RUwID
KKbbWN6QKkXERqRyjGX/CLuTkWhSierfLTjjxCTAYh4EiRXM3EmYr6wtZO0mFkSJeEdFnDSgP73V
PSNEQzRk9gnEq1w2Y/vUENnVyI2/a04tJUnQaW4rZ3me1AwKkwTAI7tGSZjoVz3CRmcNlR7k7n9H
OIHH573pohZlWwzkc2MVQXkKLAhcIa69VV6xxGCClBYlUsq8G/qqhZWN202yj94G0FY78IUlR8Rx
f4bdSo5Nsci+kFcSBFYfoaczHO3DpslrZkK+EPYddSPkq84Zd54o2ebiEHwQ3EaIMeIBdvoswRuI
KY3klvvRoJdo2pRbB0jde5YD7QWLxSV+33QoL/F7htBAWadGiFALC4Y1raJScyEgPH0faBJ4458z
/ITf/4NmLZmWdYH/d19x69wYExdQRnBNj5X1Z+7eiEeZtnnupNJED5wJy24ao4Lv2h0B4TbyPtqv
/NWJ7kYwVKsU1yHKoLoC6DnwRvga6pRVyxS1IEkhDeJyKyRRykCYhSibtiEsyl6tyYo3dGY2xkHY
Z48+rekVQxSMH5IHYuuMMH9fy6MAMgSqpyWCiqQ2Ih5/WEOSz33a9GzAe5qVZgiup6fBU4JSjjwW
z1n0lSYxifvMiLNy6peeSaU0Dn5AVCGFTktP1HTOIFHI+3N6luhNVjV/KaVLX9fd7LUHJ+71nxrB
zRfX44lFbnr0+ssQtznvZ+ep0hdPgGbd/HmACqGuxPg8/qg7VJefQ3Swq6Lu9pCdOwReT0oz3A3p
yzykuEEbdft6ND0577gE70DzH/Fbv+buNX0cDAhXd9N+qay9/itx01vCINV135KYTGVE7qDyZEFX
ju1Wfm5VlWEFhgZxV8AniDwgcaB3qMfvS6vBPDo/oHWFZSFZ3OtaQf6DYpUq+pBZDpsO1N1ttUQM
+aYEwGopdgzEKud+1Q99jISpFYkj2MBfmsMOIhsl6cKX9L4XzxI3eouZiqsWRn+RaKeBWWLLL0Pc
Gfk9anAS7mxYwVuAP7AgK+6QC2FmYVW79sX+4dCPqeEhiZzob1D/h8/Il7abTlWA0QI7asqvzfCW
3g87X+Eg40XdJ+F8pldnKF0aa/5JUnQzEON5SNXAJuSCTLyWR6N5ZbRFHs7coq01/ArxrPN9sHj2
2RKx4hc6BOHJ/5lBUs51rlxj7uI1dqcGDx6vk7LVR2j0VqV2+iHNe+isThjs2oxUMX8RhUhRuO+8
qeghMPM9RaUy447laMzURkeoLJy4Pk2JxdAMLPfEQrXbsGbHp/OOE1C0wa+JYmDGOhtgrJGqTQbv
dm0J08dIZHt7Ba6SgywTrQAwfVXxnfk3sPrrOiHE3lbQSOflGtx7dJ945fRBH9OpLvf7ojK/2e1B
QZV9/e1wHRPkWRxvIVgvvyJUHdvof6Kx2StqWtwot0zcxII2L6JdC49rjAkMytNTA7wiBitsfm4L
WYZJ3QQMmWUEDgFzRFPA5Nqz4ca8qvrXi9MTBCOw8a75ysTj22iwetcKIHNTjvO3eew7+0cLZJsR
PGmLT1qZpG1fTxFK3yUoyGI0GKjUhOYyaeYR9KrhXgy/Knw1q3Od4C+/O6P39m4qJqEtMky70Egh
MPy7CY3LWpCMefSi84wsgsnvtUgPnn0BcW6wOZ+Mb6UYXUnZ0ZjKarG5NAtEjUyC7USSj0hB1p+a
g/PTkn4srmy1gtV0Tdr5ltw6DmSnBX1bym5BZkEwgzIH3uAJbQtdz6JeMK7iDFX9okdT0WTogAOZ
+mej52STsOqTMB53hloEc1mqlun6Sos+tJmBazLedBTI5mHDKlIHOnkR1k16EPPByd8ZBTpVJHIR
MvSFE1FS17jmzwMBn01SdxwKal2OEb62heqRE72YqN3VLSaPOF2VglXWQ1mH1uSl8NuWEaaimMpc
gdvh1oHep/ozCaQ4towVKFDJQYm0SYPZ9a3iJnIYh3EKSZLnbF7v6iqnO2/JWJmobyoA2jArOXnt
ZBBDNumRL9Nl+eiw9ggz/CoGQNl1+qPlvw+laU/lMI6BFm549OkJROaPSu2RBkbQCDbKQtVFivvj
nZuSMLf/lqIUWfV3755ukpleUAZBqX8ffLABkWOFq2Mq4hlI2d6kmrwbi42ypWSZBK3QBe/RWcZC
OcCQvtuFLAZmXnSYXYDYeYV+leEEPX+nsFMnamZCiprJkP/cFjbKsyHg0B+zU0IlbkxPa+Co14p/
p1zjSYm+MhmftNBXcYTqXmC9Qrd8zu2xTax/HiVsgXnwnInqRB2r0+l2B5C9jc2uVSy0fa4bp3l+
crf7NLqvG8BEfSo+T/7/DBh6KILiInQCeh6vDeIBEE+MFnrVdCQtENXtnvsIxv7p3PtB2APfMo+3
X0GHd0BXIK4VmQL0ELPrNhiMgfwiaEcx5NnrtfCdglZuKx+juaUH4ouoBKwmOu21rJInRWxNFQf0
9Ro1KhCLed0TXjZL20aWaJ/3ofsK+ZLcMFF4cW0HSZEi/goA+E+AmYjJmwAORr4+Ez1IGb0NWujG
A2OBAhEPqzo6OPXoAMqrB541FqtblKHEzrbXbpauFonoLVUW6ZjNu52dy+cGbjnTqHCOc73BVXUu
VhmED3lvvmWB2WCDCu781nc//Oo4/BFjM4B0q8wqrNuUXKxrroTs/uHzYKObyuVz7gSIP9RrQ29t
I0Lc2FQ5Ox1KzeUdGNLamC2VQmXYfl/S2VtQD0ZQOYx//GZzYudmGreEbBEMF4evu3hcoBxaUa8p
zdYNVZMnkYjxKJlpbuyLQpW6OzBNJNkZ/u9EBxS+HCycKERQ8USlFEf3gXa0y4XKdxg88GKaIIoB
+OBB0dfEvtCnHclXei0hyyvPt6NJlSMAlT9DJxke6VNJEuOp9vnLQUmtX1NnIRJu/BhIKH4T4+m1
Bos9Z1YcgpU0WuT70rPWR0jUkk3kNt+eQDWwt6hNtua/j9greUQRkamTkHT/7bG6xGwxkp+QZFf+
yZsWtZ9birBaNfcYNG3PRIu3vrkcKsJVGTQvD37QOlfMsyuOPlK7Y4Ao06kJDjgpoDqULhz+kCts
jLOfebodjc+ZUldeBzR9bQ4fXGFM9+dSq7iVUTIIN5Yn1lBWcl/SeVJl5OfgHZCAsZVb8yylT2ED
C0wP3db2JeRhUhjHfJ5N4qfq7E3las/dscxACPxTbFNbl8M2n7oIaqcYIu13VdBANjA+hW+qgO8P
fTuryJvHpsf/IuyfXFa4Xmcxyk3sEa6CP5ZX+6qatA5xdk2PZRYhESTalmebTrIG8yOJmlGbLlaE
wKarsXMdrLsy2IelP+Xi3urQBqXLpv7v4XhWmBY0AJkim+FcNuT9TRLXgOl1KRVAqx9LNR7jv1dW
pUzQ9XYMCb7S8lqVIofi1hd1i7aGeqxeKuCSneHNRTZQ3jB1QSDmZMEnNH/bwghP+TnUnmVmbLuQ
I8NMRF6OQou6tbPi9QhGWGHQehwX8iJt+GRhazO0FhmdpGRNXMx6+m4tpqHePmeKBpDA6lsG4g7M
iVuoxM7x+jYHWQltF1iUXwjUXv+hmeYmSvIsn/x7DcPHiqnLsGMjQOvfvfQO6t9hG93P9JpN44Ff
mnr9EhwbZZAd38tmvW7wGkK9jcoEQ6+oXZ1zYwICsN45VQRsDocmLxN4Mo8P5cP73GsgKakxygqv
NMqs+YiA7nMKHQGwx2BULwEubiyceEtdDSoDlHRSH+7NhsxLnoeN71L0jQNRp8ALgqrYUHoddiI/
CMEEgPceAtrAvqsIhu7UQ7xj601RIGIrxgEkY2G0uhgitfXVj3/prC4yJNzj9dqQuKYn++xHrDCl
LJFoIA+cF/JBAo0hLEgJUsLQ1dYcWtzP9J6YZTQ6mkifc2WXFR+BrkHDSh+kFMHd5RPIvhZhXC8E
N8dh6niqk7JOyvOY239b6VbD20BAd63Oh1qvfLzxJwgxR6tF9V7Y6WWo+6MTUdlmrAnQ+mNumoyQ
NcpR874taVwQ8rN2jjCISNCXR2btYd6VEnBuMvGifHJWclMNGGzGgr/1M9pGGYIgtH/CGStWJXgm
h2VqY23zgdaVHoCV6jbU0a4UAZ3G40hv4Oje5RG1zhvCXNjrCVrVgCY3titjRikauooX4oaxTbbY
zlaAmr2/55kRa5sFdOAWBVzM6QIzHn5rom3UkK+sjkneZE+c75fZzu9TKJgJyZQ/Sh+ct+X1BbM9
IHhWMluNiZGMNEJVV+LyAEoYPjd3GrvGcZytCy4bVoGghSeAwQklzjtlSSBgkvWspAP82Xf1nh64
v6n7TFNZxG6AUeI5YNn2JoNoqIZBIoxkvFK5pF+0tnG8CfvTAWB/K0ApiMYD6XzuQsT/rOXn87al
upIzaMryHIXyfOVAsoNsJxz6tORPv9HTQtBGf+bMeKOnKlC2GuwcwTvds1E9CGC3sFtkRkOaLYVA
HakE4uvx++x4DVYWDxUAdUtqpNPcv2uO7OA6aHY6q6fQCbKCzDEgSnxoN/pfQLgLk4lMEe4PKeqG
kxpwcHaO7MmAtpJtmiRiuyIK6t9D7mVXUX6JtI5iWQZc21ldk6e+3ZmBBp7VnX3pyKMl4x/IeP9/
3mv9ZOUk9j8JhkfZEXPXakVXCg6Oc7nOHXNeBKR9NXvs8e6dmvf6Z+0eA1CielUwUvAKwfq5GRw5
JyPnHTRsi9I06/22sNZaQjRCHFLj5av4wGBgwgpHHyR+xTJuDJHJsuwikz1xfOnX9a+CGfhdzjEZ
V4AGOZZCGNN2RwW4KjCFP87lhpCjFZurf+YRXSLpvwS6+zXSO0a4cWAtcHoAm/8Upco7nzjqfXH+
rUxj/31FR7bezG3CHtFwYyNzYUWdd509mbX18wOQMZ8gJIuyKZrGyGqK79/+Fj9x5zx7RGNdCCMN
ceD0ylMnntkR8uiGMFY6bY4bs4nuC6TuE2gxxXiU4BsD1Hed4LesT0QdulibHnn4rJ+h2h6wueNa
nhzSeWz4MRTeRGgXSRLmLhDrqZ6Brej1+wT+c/3fDVDT4GnjZT0i79IxqIZS73AZa/V35L7LkYoY
2sqvtoTr3E0kwywRajzGGqK/5tCv6ib8VLSt3epJ5ThgIhUn96GKdEarfmJfPR0vK2VK6jK+wH8D
ieUeU7MSstgM+HLqzoSybFEd8t6Yv9TzSY/81CqsHiC+tJuLaKp/mwEzwT+dsnDK8UYYIifnluHv
LXwBP9N8jKDgTu2k7/L5rTpsYLZhd7zPCpx87+pfZSUfq6HsSFvYzZpCm0SOVEnX0OyA+GFm6DEY
GmdwwQHrybz6U7uU77QxVEVn6jZhdL8/ebat/RtHr4wDhD1V7ghX3dgrZU2M4TCbwaSgu/t5GW81
MtCwEv4lc8fg02FVOQddEGg8DxAF/LPotQ3YjrWl03YltxJJN4q3NQzyRz82fZPrbrPLvXHNjsmi
Wy/C0Xo8+4KSLVKh9TvkfA7iPBQPvNpCFmhWsCHZuVJWCZksiEfaBy0tcJOcIqBlLrvINGjnlKmJ
YO23wwcacKNSNMLPviEW0pRuAsNFZUzpbhnIZuQcQ2M57iL4w0h1HhXPgtFsadjL7rUFuRnzw0Gr
KUIOxeiqN+koP5VtlAEfjlxVvizzZNLiETeSUF+p/16XLB8Ev5wEGwfBFv5OKUw38JzgJqOCydE7
H2ZPzPfQhsm/7v0FP8W6vYhslDoAv5mtP2UrjcuSGKDNz6Ef8z/vteIjdG6mm/a8m4/zWgqDv1IF
eF4eKpgCYWBbrVU9BgG+/Rr1LqIxxehqpgLHUaVViyAGSfbgu2eK+8Z0aG+LqfBeOuG4wC7xkjhK
LrrUO+IkqjFPhr05xGjM3ui/74NO+JypzcZEo1NHG/gVD1zWPveIVSHZXpssC0tBQhgfl9gqYxrb
swXsCDygryGpruob+mQyfHD4OXrkB+n9Zg0Dsigc6kVwjTPf8t9gaf1J8MZFAPCOklEwRiLjOID9
27YRD2IvnM9DjTOoibHXr94wzRK1l0GZGeg80N6xRBj44YWEHXUh60l+io7PLmhflsUZsqWcrS1f
bpbTkOtCIAraawznWRyLQyi3QdkQwmT7BExeovwSWog5FxLvdryzbk6r5CtRwkYMUrzqM6j+DvVP
QUJEW+OcvG5OhP3EJxKhn47TaKc1yVWktttdnc6LMJeByJa2Z0jc0+XgztDbvrgFhL8H/rg6vXvq
80ip19d0XddDaJYqdePnYkhYiAQI/RA84jGNQJ/qc7S4fo+2OftSDv068cxkwBG2W//hkDCivGHe
ihIPPp3q+VkOvid233zbuaBhJMv4QQDdZVNJAEnPai93xluEJHhbQmPIrUqU2mdCtydRA+1D9DFw
FpPDVZstOYdckfTkyw6DNgmuSEhjjavYZHERIZA3ccEW1P4+3XC9++cdsC0JmdDt7NGFPbk2H73h
ZmpTar5Ja0mrXhblK2U93hxbz3di01oo7bQh0eItHxh4SKS6JDHcWJbf55US+df9sYwjP4f5gxGi
GHRKe7lucjbbPi67NCkNlXarU15ylacBKAWXLK4dFJxXSKmcviNMgvKxZSdXxdT2HICahHklLuEP
h+wbvJvn1N97MUTmnqcru7opBx0zo9ah8SGGPwCy1Hef+U0wiwwF1BWzMQjB/5d/GcD+1JyHnc7i
neKzcrSS/hFr8Teo0wdcpdNkuksvUFXdteJCA9V98faXSyugNRM7soPCRItAcUPSc+K5TommrPmi
KraMK8cqqtbtNzEp/Xll/pqC4oN+qfsD9HlWSWNgSjZhS/f+end8DuUtH06X3HR8lveYvU0VddDb
8dW6sDOLYQ/C3iPlfL3EeavKbIyPep5WtTdoCj0L2qH+W1A8HqGWk2+nfkiOpzH8652PS9ytP8KO
V2b/8+aax+INVJSJqDtws90xKB/6FEruMC3n2AGG9iSiCaEUwIe6uiZFDW/0W1mJOKVEtoAEyofT
iZY1HwtpnqJ/07Go5hPhv17zstenPV2PrkxmLmFU3tJkG4Jdwd1KGWdT7Uyk/Er2zzQo5zny3FGi
ooaNyKacvNOiec1dlwCkLobnf/WfVU1rmbYVi1u3uz6+lNslLjbfCdYV6oWbDeNqUyuVFHmN6ybq
3AZrT9RNkfMvLCT+QkcZmKDiUUoXciE5IbDXZY7w+Jh3+ZVtmB3IPJ2s9jxUIwRLK0KUC+xs+N92
JMOUbovLWkOr01gGIfoDAUezBeKraExauWCroRILIEb4aic+dGiCXUq9ZIgSmbHDZd9/mFJDUKfS
XmgFQFvFT5ffU5lwjCiKhfcooASaoINXl/i2nGac680AP5inBfgwRcCx7eMxLudx4rEgdee+lQBH
zSUhzUFCeVVW1BTC0dHdWHll88Vb8Rt1VOGyFM64YF6loI0W5qgRkRPkOgzK4sCRecrkIoNyqGz6
bb4lNE2uIqoK6nKWbpxL06sgsEEBlsGkODL+ou88axHrBSvge3ZVScLDhi881aoOiyvbjSdPE3ZQ
lGY4Ss1rd07O5Vfy/PyxvKVtM5NCrgtJflvFCyLa2wmBe6rJS4CF2JVDrrY3gSjmZaTr+n2FCmV+
s8xeTUfyObgDtc88DHcdYP8K1zi+ZpG9J9rp55pxL9igg3gCU2/wdwC3Hs8GUmu5gM2tKYbru+Ip
y4+YPGIw6OGSZqbscFzSu5bbhY4e0Uec1rFZ9oBUW6a5CnltvJ7zegdPvk9JEdTwg3gtQ7q/eI1l
o4ZQudex2kO5FGsJv3XksRHkMPp/NXlourpWFj/NVBVHSsh1ZQZhUUWsiXvZugc8fx7hRlheBZqr
zLuh095+Jgo54U52WIIDkawoYeLkBOGo/7dj07zKih5J2acvOYJk4ba9C6336F1rrXhb1csQ/dVI
KocVq452Ek0h6w1dSwjK4ZaoCl/vbpkR21RQb9EveULZto1ABnv9UZ70dptJP1b7usuKcTKwtgTy
VERXFuoja9dHMFutXZNa9YUnJTv4WmBHX3r6HCS2UKMyu7UkRhGiePJMMSM9eWzM4stI8k7sz5vn
M/h75picNeV4G8FJts4vQkdhu4f8+IpIoVGrSHKOaxqJJWicZEqFNAD0Jn0i2F/m283DT0BKBa0V
Xj95pB0vZrhwu7CJYoYPHXG6CN55KetipGAAL29FiFnCr1oZCMqEMrkNerqzHkmhGlODnQCWOsPX
XdcTjt1hQd/NjbS6hXnBZPuqdJ3IuqjvWejiTOIgrxH4+nrQnenyc0FjCFgvy+TUHjHA3LFvg2Yw
250dusp0XOJrMohiDxytE0a6MMwcOqynoVoLNLr6796yut/fzuElyB72exhOZb8QvL+Yz2tUFOWf
DUssx9yIIRS7QsLa5/FEv6kKgZUiPi+TJaVTVvxXXo0kigcGNB81YUqbyD2Kp7LneulrNvRDZ5Z6
28faiNHfWY0x+tqZ7GJUhlKhGE60BjGFUIAnAxJ/4HEV3VSKHjqPTD4aNeu5DrYYeifww55oyujb
mgIrRu2nzuSv4qWvMV7LAaOoT1lykl4yh3FnesAzfLxMfpDdo6btJHVzfo5k1owkM62CL6P7YhaI
oEad440IFcE6dFFgFJnzZWz3iU2IZ4WmLa/14ETfi6mzo8IPjAZNpqZC9VfLa1YkGNIrsAbmTy6p
z+Dun80CRd+Uiwj+G2xMEHFVQ2u9ltRloiDVPTZ34G2TAIDNmGKEy1n7G7Pzb5pPYjbs3ymygkaC
slGgz7VeOGC6HPqsbq2B/xmJAGtWqLQQppQEXlgmAN4tRtYcGp4r+FmZjtlGinWucYFA2YfJ6ceo
h3u3CmEJadoDCkyGW6XvxXjRTLPfLp3qmvsR1t+Cv7W1MH5mQDryOlwc47whg0RGA0G3e2EVmVNN
iowTmWcofwF0+SHcxeZCazEd75Id2bvPQpmJJj/46uJmVjfGEWOV9SgCOxazZr/KVHrFpFqEd7IK
aAUm+kACMe9k+b/DMSYrji8nK7J0CBskKpdoTOv5WCCEcPrJt9FR81RqQZyfSmcfMaNTiHcJgTBa
TgzMtkyigE4NAParo/OgLqUx39W2SE1+SgmKm1R9Bl25G4y7BodFecXsZUsdE44FqtnbMgPZ0OJ3
uFIcr8RZ3zWXrb4dKgjSzhfCEeY+lvHFYpPX11iIwm1CmKq88oDRhq3RnWfTPruSedotj78zvrx2
9huwW8CbVXCXzICp2PDxypZ/semCZ6qGXXTogAfkDWLRbj0hjtgL36O49n5SBtjO1+LjsQ9pU6ap
G0gG5aUutRJFaG9MhUw3nUG9832VWAFoNr87X8gmQDgVylv1deTY4Iz21Bo9lw368u5rQKB/i9OM
AsuIPGNwPj1A/AKmUN+uvEYxyZ3UC1vzVUTx1t+xUDgHa3mI54qXN0NxU0fNn1Mi5A3ydWKI2Ic0
EbNT1mFyv8H+dwvINUBet7ssK6GbcFMDp6bKq3O2EiEgXFPs66U8P/B6S6MmYu2FxyTRUOAi2hhX
N3jSaJUgmhlO0dOz53H2OthemP8U8s9YyZLozgysVilpMpFai0YEHdnSZzxPhgu43l7agqWSJ2Rs
0XJMzsa6icYW87yqEGnD5205VqRo19mFHY3ylaLBDlgs4tvK1e+j0KEj4n7Q88Cam+LfIppKsoz3
ulQUGLKFRKJUnyf+3w547VqlQCcyn5EM5o8VZ3FTB0+2Id6umJUUap2l9mlWIfpCwbzi09Wrjr0X
9qKKbgvlU0gWfzUzasPNI8AHEaC5bBVimSSVvQtBSlMq/ADMSEX0psCs06A22q0qxytacfwTzi8s
DPnNL8LxmRrwUTVS4kHKhj1cr0YAP9IjE1+MFbDh9dxdSfr3Jag9VG1jCBuhGM5jVshKA1D2JebR
Zj/Z7nSe9w6/FdVM9xmQzYTMbD19eliUPKeFOclmXhMWnyyFxqVkE/0cG4oWFAW+omRn3IdgAoD2
IuDpaRjzq2NPhbgv63rSuJsBnTcg5O2KAjDwA5UB7NokGwrtp2sjairyIHcDJNAP7YikLTGcpctQ
9rOi/C/WSRAPbJYTrdQ1yujePK8S3Ps23K3zIKx6Khr9qoUsdKrkhU6VrP4AuFrf3v8m8423gFLL
i/QuOCgjva7AHP0RelWDMnfi9nErxoz4TYh7ST4yE6pxPUSWSQz/f7Q2RHGIySnj5Aer0YzDVEkD
g5QKlFlMYw1V/x0A+gwLOdOcWBlHKx9qDx//A8OthL33EKsy4CAVUN1xyl9jviKP9rlHcxQLYL1Y
vjZiIm0eWc+LQk7ZaocwC62wRL0FMa8kZPC8NEB2Tg7RRXm1H3fCf2tPtn1BmWHTIzpkovisuwnJ
GdJTKjBv5pPQIFk406W6XTDZtSNvaRwGdPWWoRN2X1J6DyVJp9Rthh45Mk+Z7TG4AG7nbeVvGQWY
6GG2jIgGj6vFjvppeWigKLUkDeZP57xNxw8LtnvA1D//eeJRYzl+eF/OBE2fDRyT1PZtXC5hQe/y
PIlerEl8VhWIGe+kk1pitWkmW3VOA714/HZKtEP1jkUttDP3hAh3k9aykPPTedj6Oh6VYUQA4klp
Oi1gfka9INPtAAS7nWWLIR3El1nSYJq8i7pieXpnlLKAE5rJTjisoOnGyQAhYcoRZGsMGT431wN5
K4kiS5+vtIXv04unA557l2gXpPQpKEIveeXMxBqTeX6cPT2zsYC9cE5NR+cBCEY6rRSxMIXZ9hAr
MpTzENTDeluZXekthqcoA/Yxdh1UUY8/LMlpiyZbDUgqf/2gbvHnnDARIIZyrmKyGLg8eQeCV0BC
817PlB/bUBPB1jFTSl0/DUH3FctXpiyERPLl3lQc+SlV9UBImmEYVb9qa+hPEQKTQYNYj/Ap7ItF
xSDnuSmauw8RiQYg7S6HxLCUYha33VpfWmoc+lA9YmL5ckRzHCvKf/DmBxVRveuAmKds6U4Tijmm
PVu+yDZcIIYfHxDVlfrS7CXe9H0WQV+lmYRqge9kJ/OLdH+vkyiSCTjr3mtE+FTk0tVJN0Oso6Vh
Vv54R/ppMDc8B0m2c8KztZ809CQyBMH//CoCunm6g7F6L8xY44jnEV8Q32N+rhsr/9u4pkx7DCbx
gEQIwufDVxX6+RXWhoPHnu+84zkC+t5IhxEwdqaW2C+lL6yua8w51HPKiC2ABYmDoa8a1XxfCFd5
Rhdh3KCu5jx3uyxWgvS59q/QD1KhIYDZ60O5gHwBnILssz6Dt81Px33i42QHnq9ctoR3/jw+SFyC
LV/1t4GQBI/8zKUmylXCRicyGk3+ynEPMlaRSkzR5EEtHRV/wNVxnjeCq5bOu9WObmQCqYd50F2f
iPZDrSgEijvq7DaxGX9F2GZbB5/OvAZ2V3Ezajnl9yIevioUdW7oUWcf7uJyuosk+RKiSDWLbofD
eqpeJEgKqQO+tjLlD0HOUGQE9Gw9xa94jpU37LpMYVugHExOJG6zkkkmsLt10uI1QNL07goPGIRr
SaMSH/qjpam7FkMCpHkKu/RHjoSW4gnWQ7ulwhIJpxuVxQgrtUkdXsNsuCVz/OWPg8fVp6indg8B
pbpQ+nhotBotCLuJxk8RrWoRbEVXNJr+4XQGvgsCsgkN/cLTvf/plZTheZHry2sWGxvqfO0YnUHe
MBf21jOdLxgufLxLFlHQea6NO9dP34uXGkdRwPNTeZ4hSKS4F4LeM5tpAI/jvp0cK1ULhA4keO2i
tKGLF7oi3d9VpKI9wx8PRKP+ODgaALQvofwBfng819VH7jCHEMbe+dA/Vx5V1mjUXRNtysK3Dnuq
Swu+pvy6Kpw/cnmSQs0g+Fs4cm12XUOOUyXf5ONgJ1uVYLOlGxsDsHQfWXzJ0VMRSMW3cP9pM1IH
iEnFflpV2ZuDe8HDTIHorxrQHSLtl/zlxiZgBKnu48MmEQanETDsfQhvPedeFQXTXb2OxqllJvCK
wIR/WobOjLXSdp1LXcRyDRAJT7oTDBL+siT2G14juSLh5BxB2GfwoyHZ9+Bc3JygsHkcAp9IUpY8
yyMvrYLbZUf4LKOZxnkMudx52HxCDAxBxZhLd2nC3uM3NwY5amXAhBcZwRSQxqULSErsXpputzo8
3hWVGuq6ffL2BKIWBFJ12o5WsQGxVtIcRNTAIeMRgLEMK4AG4k8l2UuTt2Gun/rIwaqwRg8bgKuN
rIE8OKzrA5hkxC0ueI4AB7kH9yMOafZlf+h6fFsHFxQkoYmpxu4CuvusfSm/tlKNGQuEm02eBFud
xXF4NHxRlAeLs6q8QdORINPfRSf5QdOy5jW1ap2JNX2RsKeLEQCTpZNxdtvPYTdCSFdZFij9b+Bt
Bbs1EL7R4OrII+o3pMbwlsJXTBVKczHXvZbCKkpi+VKHIe6Pkt3IE/1/BzxC2GIGOWSCyZTQvij/
b/xdXJEgvjU2vGfNzVApIh9jSjN2FofVi5oR+xwUWGu+/Rb+u8cVEVGnAcGYcvV5BsdI1KFJZnFv
XpDlS6LY0ct30VC0zk1E4iHjUmJJE8t6QtEOEClT6ZGBBWoy0ZzM1eBcstgDSe0iSgD4rf/s8lGG
Ulpcur5tcCuyW/tdRqzpCj2P/c2au31VYQorjb3pw2j5Ob+JmqzN6PSsYdtqmn/YL+lvpiqubOl5
ULLdmVl54k6hxEBpL4t2bIiSiYpnszA4p7MxPRvd3ZpDLuEM5FkX5nI5MIVgqaQu9GM0E2oe+e50
kYWyRWHx7W8NJMCoIKlBxXTxmkKqq/TULEQ4+QL5JLV73TSo6LAbrSrRYjYBaoWifh1Dm5sKN270
Zs74y4rrViNTF55S6vmf9sFpt1Ays920KV/SbhFpzGXX6HYAv0au+LMuYlibuNb/yVpsAcB+7DR9
iwiFUO0HNMDgwuruhcLQEmxbH41PcXseU1Hwo2Ftf6Ybx8Zu1lIr1dThNSjghF2V2cqX/G5SGOoJ
oOls8/IbanpAWBVbVXUxEa5Qojo9Ln6PDW62zFuz3fGDVJjPIO/0I5UEVGkuWY6rLYAe9F9eT53n
EQkWgKZOYb/Q7SamDL2pv3LlspkIgYID0oGZ7Ww/i4iymCpMXYudRFrSkjq//UONjH2+WY8Yk5XH
Mo7gaij5A1uZBg0RlJLYiDAU/lfVYqRII0giFe0RgrtvbhBCJ/J8ow2wQu8ULldS601h08eNyw9w
QRtWT6FaAfzhDSmpKH8YUQcsaZOSLkTlvNcrbRLASeDCqnDlH1Fy54arhmfoNjJEOfDawIg6E1tq
m30WooItO4oLL4VUKIaGpzqsgza1gF3MpAFtd56dOdUqiERldxzBqzIHh6dxxOBVpjsqyGs/L83u
LGlIHq8YCzmzAUpHAFmUETvmdd0KQ58xtVBJUmAsCByqPohX5D9JVzyUlrfYwh2N1sM/bDhvfByr
vfkTq82bMDgiK3tIuUcIWF/pgDXTQMK191eEFzM+cJ0a6m8srC7TCzbWjYBcobHZF0zE/RciJbKq
GTe1ipBB4zeUzQjzcCmChdlmX3u69/FwW7AQkrWqTOs25mXNefwVOMUBk3yYp/bPI4I4LQBVcf6Y
G6PkHhxXbzUwlRBt2YwlpOfu+JX3wNgSt80aXzTyBpeGH0dNukLgAA6p9/J5Cl3DhKkB6/QxR0/E
5DxymEdifPdyIy6YFl64lk8+tj0swUtWoXKZQevzYCshMBG3G4VJ/0JrUpEmBXjk/NXrMt4cLtp2
aRXzVyzaffygMKOvqiPkRjlvO+Rha19VAOJhqWizBm5j5wqB/Az9f1lVKeDZRFcn9v032KqUhCx/
xkCRkqipL1cwt1gV56Mxp3dcANZDrhyz57GgcjrYuxUzAdYWq5Dw7W/FSgXcj/058cO01KAtLrf3
ikRBARnTcLJQh4AZTWKsWGuhaeK+io59UabTE3PVY2BCgz12ynBEK8OSzMj3hvpvKxMe9nSazMRx
xv8nBGsW2bXCQMDU5E9RR/eVHCVUcpnNARDe6Hv3CRaVYHnUtNwJ76y9sJbw5hTV8c82QbkqzAOx
i5iNhTInXyFCU9RFhbgoVunHSYqNGbcCyCQY1sOjfnxEgp/SFc3SjdnxkjXbeVaA4b6nY5mUkEBV
e4LbQYPSq9ezoRSFqmDRXeMbzEcM0jvvT3fGHcw4Y8Ht087VN6lefrdkBaH82Va5baKebkNvW9FQ
x4k8N2kzyEO+7g1OzTfW6UBgbIGNUxAoSigltUR/EunOZ9miGd/v4N4gK9rDwzktYORMzvFw1ov1
9Xl4PHZmyvcfRvpf1tw/uHrArnr8YsiM1Nny+U1e5GIZEjc93xIiq5fiqBAOnaPROIla7T/5Utp5
LSx6evz1tOGFDV4mSR3TD7zKTQUcLW149qEjcGMMHeNnTz8BYxmAY7ifmXJ5dDE9ac70rei0l7E/
X/zG3zK9vtM+qD1IXHNfGjfSUCodUO9VkLpUSlVetK80Z+N9KDCjJAbhSMib1CATlCGHUmBaSWhp
G6MlfpDvEGnXnbH5ZHQyzs+QoQeGimGzPzcd4kWtZS8kQLlyoiSCSddvdqH4UnGX+ev4yc15A8C/
BlDeUaqD5dzdSm3WypsbURDgCMfRtdk/qZWOX96M09gl/w0yS0f9zuAJYEl/n84XD3BCNM6aqse6
vHxA6Ct4eTI0i0w9650cyuzCPLHJ/1bLhHtV8gsdapoQZpj3cwVN0K2094WA2dzF19vFVE9wB0Pv
xvpDVpxZFUDqkCOoZ8VhUGrrEOnVDnaJhXnmPr6JaSvNO8xiKVEoRSZuhT64jbOj6n9n9vFeH/nr
mu3u8OYgJ7D7gkq7H8HN2EIPM7Hni2BfBg+ySxUKKuJaTLwx/C1JTKVM3tOGt32kbgl+v1uAM2av
Gw8RF/fAAiM0hP744z+WyvuecZomSibtx4ipGGetZqA8nXwgem2InZGGeR3T0JZ68H28ztkMwBdR
/XeOAMGj8XrCQtRv6w7FWSvqRB6h/M8MziXUGjcd+RvVXQcBEyHtyv4G6yNrLkTzYfFMF13naV/C
Bwiu+uZSKimEZXJs/Fp3jWJ5b0lyCYXNvU0aJvXa+pw3ypJZz964sU4JPSTqozAeqodQxWljJhY7
2daQJs4kY7YqmH2b6LDEGASDuFJ3VjpmGVciNXtLX7V0vp6e5HRw82KRt+mnEQoML8sB283UHzOW
qyuBsLChmtBrpYsJspbG2H8h0JIdH8VDAsscOFnAu1a+8xMpbGecInl0gUkB74ZdQDpHdUjoXKrK
ZHcykQyMZyRoYzx4KDCEqKVElkwy3f0VAL6j/uWxMiRPustcgG5slx5GXvi2NvgH+v7o127N7Csf
z5ULN99TZgDe1mCPykH4U9ciI6ssF+Oirf9v3AijcyjZii8z85amD3YhU0oPNVLdZW5o80iV7haN
65caQK/oYCyKYUzzND4ZuhJXa+mOnMu0lmdyXmkjEPwLJTnbKSDUTSGvTsVf/WnEzx7lO4QwxL7c
NSya0pGrRtyBsHGAwOfBMn50Wuqd2nwHfhw3lMwM3xXJe5PdI4eJemj80f8isbl7Xn5m+Ej8tIGM
OxS9t1u8DGjIuI7pga3mBRyZVwVkdRNrADWdu3sMpnqxwhkBsEwf2t3ns4ssF0oYkRrckugV3TFT
FF3fwfg7iupwhiAMO4AkAW1+VUwdfkgATAAAxnmuWgSKDzqLt+wg1Po07kFIQl5Diw/vgjoZKcl7
tJxuz8BU0LbPQaCrhTS/YGlUyD6/D8H+SIHxIk0c2B+B9x1YL5sBBjepzthAjbImVJHv91OnBnAL
a00e4iYNucgjHf8ZJU561WaM685gg6ciSadUFjqeWeMTvNMrdE55I0Nd890eWLgw2vi1gpkvbU/M
LZL5kG8lUXCZNQHR0xRk49PnU/Bdmd0hU/3d1R+B/Ofs8AraysFysn26ideoBiMBsiylkNlG70oC
3jUb5M6cM1dU6Wf2eXDU3G/ABpqKwrzscq6W8BZYl3Fj19umNt2JfDfHRgFUOt1Ti5DWhc/H0vtQ
Bqyu3CGEgL2GOCqIvU7TyltICgYTos+3Dg14jl9XiS84uCKn4IAedI7Pwoi1CtXKSPf3ykJO0jEv
LVMzdpIqF2uHQ6SzvkWfxDsgggzX8F3+f4iwW/hfOuY6I3lTPr82hnLGnxlxf0nOrnsKUUXeNStC
2rQ+qw8U8ZKhK6TcC8Fy14u5sLmEq2rL/g7lo/eYtGdhmkHJujcqrte7Jkkc1IRinv2JrkDYZf5/
g3LuQtfWoHYt5d5ORF4pKuih/N+IA8BNUld1Dw86o2MkRbAjiVKJWLSP3zz6Z31Ftuu7BSOrDY1m
7U9IdSzpkm0kS1VfYMLu75JCdKPRaMEOA0DCdAPPxVl8D5LkenEMMwmFUaPZSY22FYIJ5N2OwOWt
VY7BNDkb9oBC7826GW1LdlI87OaEjoh6NxtGV0lnBgMwkEZ+xe1/FtDtiixc3RgSWxaQZS31t6UF
B29ZQmeEfH4TY2BLOfAoNZVK8oV01hVws77jt9TV01+ueQmuEJrAGtR8HoKiTqolrBhQLT5KQ8Cr
ZfkRwg2j/23Pu+zbP7eQ+JrjUZhNWGNbrzmFaErqyE/LmbmCjFJ8U+kMdd7DNSuK5/BVfx24670T
OcCjNbgmF1G05O625m6jcQLt+3ZJSuKeuJTfPek05ul6i4s3J8r6V/KpF/UYn/WYC1hhJLmiuBd3
bzSJdBcpjQlGCIb+Ua0eqPPECK0DFmosRwfunxIIsvMnhJXe0wr4zhCr53Rcf4wc/1tgjLOMZvOQ
MtGgG1NxJC0xTnFnqilXqlNw/K7pKv/GhvJvwDJ+mr2P0koitbWCHAyLJ9q79+YuDbtGLwFHUe8V
w+LF33yW+0KZY8yUW/qF5Sbj9pzKo42WwrtDOGINz7Y17hDTxc8H5lI+aolR5Rvx/lc73/HfXRbm
zYZKE3kDVQ48318b8wSrAxL6t+/y1HceCzHjKIIa4xFOJ+O3F5J5CegfbhwCBeKZSlLagFkqwiP8
QcN2N8rNq65J5/zr25QCzHh1okIRCABeBdqOMcei7ytWceUizjS2ENXBKcv50DsEkG/GtpfxnXuI
PukrjagF9/WytAMgaipThX6BddWIeUqgw2jY5d2Iukd+oeEDcZPOtbJrKf/chGzw0PhTHSqVGMOd
A5sQ2b0kAg5bPq7lPL6uaUQqXUmqYMUOX8XyISz50ZXYoiLIY4OUHBwI21lGiYEHvPKOnReFGDsl
bjBhUJ0hwqhYYY8MGC/jZpFOEUqnIfcyhAZYNVfdo4NtuPUNxzYzLl/6nmGHTZSeuCkBjCeLyQcY
9JhPlLNxf62bhqR8hXXNqCCFOhB55+9x0TMOeUqXkuVHXZjWNwXe7PrroBAKV5VmykjEDLcRhdpm
3w2jsGlOBn4fdq2zFaHemCqmJYYDkb8f8lh2RpOb65bHeP7nTz8A78bUeEHKhC1L5CWwl3/OPlp1
lnPTLkCY4hmXp2+DTuH3Nd5ZTb4z8yHUHJL65DpG1tjdZ1q8XY+KYVV9u+FBe4AZqVN8WV1Q3pxQ
7hG1P+0dfOAWKWf1sHUyOYs4Nreg7VKXuIrb4ToqwtgKQNtAk0KTGJdGMmS3aVv9Tq8dVakpLADm
3EmIIXMpMDN2UFnc+cRownPDUcsSxa35PJrWFHHv960EwftFa3jGoRnKjUWkNz6eXoSDa2S43lP0
s145wWWuv9upB81MRWSr6OpcgsgodujD6hzqmhIKguZQf6zMKdNy6onUgJ/dnSBuEN0imC8rMp6m
+gpVkwdTxM3Nul8jovY5rrUUMU7cxgW8sFEh0F41vZzfbTVBty+HUmiV9APxHduevFPVL9fvl5Dd
mQCknxHp1+JPrxCbXAWmayWaiTeg6w+zKtcOesZ1qrfbCS2XqKI8ZaZpnywWYya+T/VE9gz3QzVp
xjV5h5+0BM+bKgIUVuX3oKtIMO6J6LPUzFINNbWH8Zl7yUair2f09qZ3FsaOd4BD2qIq2Kx+fXDA
P5e6Czw4HSnbgEzgFRerLCR6Xpy0Cxmiz8MIAcD/PoEAslB7rgV0YEtb5jSQUm4P/Y1qIBxxZFlr
Z//IRdWDolZxU+uQdhwPFaEG10i5UnaDdHUs5TQ8J0Kyo5TO2ilpcTky2JwCZP3Lm9zA6sKAODOC
IMWHULoBQoJb+iWcfB9Wf2hbDIThuyJQqXlIk0crjUtzleajYx+g3N5rcy84/DFFRdxdwXwadlGl
S7N8Ek6UzOFdjpMuAwsiUYzAEDNOzNOwXW53XgNH4SFUk4Yi6Y3ck06egEuhaUY4FMgPsoi0owvu
yHcXsTndLjYPxOtgdJPHNJoXDfX3Ozr3nP8KU6o81W0EWtXEDdXylyuqVgDa8C14tcsW7VGKL6rG
qtSZNxuk0L7MRk+P6ZvdnEnEpwMfFwYMg2q2oLSfoqJWOgIdPnDIYLfi+8UgheBvtUq6bWND3uo2
pZ2hgNcrtB8g71gmXTyNZ/ZSL5Iud8BOTr8B1k2Ijk7DxEIQJ4Wk7L2fPxTIBHbZenZ9ooYSnl0N
J2tb7DNMTUrDz5Psf117ef4MoY6wwIVwota3UCb8OO+PjC2QGV6oIpv5vNsR0BEfdsEjnM/IRpVX
p4uvEkCE2bj6bKauv7J1MqOYYzre
`protect end_protected
